//
// from command: eteak -v --gates --test-protocol -n poly.teak -o poly
//
// Generated on: Fri Apr 15 23:03:34 PDT 2016
//


`timescale 1ns/1ps

// tko0m32_1nm32b1 TeakO [
//     (1,TeakOConstant 32 1)] [One 0,One 32]
module tko0m32_1nm32b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  BUFF I12 (o_0r0[11:11], i_0r);
  BUFF I13 (o_0r0[12:12], i_0r);
  BUFF I14 (o_0r0[13:13], i_0r);
  BUFF I15 (o_0r0[14:14], i_0r);
  BUFF I16 (o_0r0[15:15], i_0r);
  BUFF I17 (o_0r0[16:16], i_0r);
  BUFF I18 (o_0r0[17:17], i_0r);
  BUFF I19 (o_0r0[18:18], i_0r);
  BUFF I20 (o_0r0[19:19], i_0r);
  BUFF I21 (o_0r0[20:20], i_0r);
  BUFF I22 (o_0r0[21:21], i_0r);
  BUFF I23 (o_0r0[22:22], i_0r);
  BUFF I24 (o_0r0[23:23], i_0r);
  BUFF I25 (o_0r0[24:24], i_0r);
  BUFF I26 (o_0r0[25:25], i_0r);
  BUFF I27 (o_0r0[26:26], i_0r);
  BUFF I28 (o_0r0[27:27], i_0r);
  BUFF I29 (o_0r0[28:28], i_0r);
  BUFF I30 (o_0r0[29:29], i_0r);
  BUFF I31 (o_0r0[30:30], i_0r);
  BUFF I32 (o_0r0[31:31], i_0r);
  GND I33 (o_0r1[1:1]);
  GND I34 (o_0r1[2:2]);
  GND I35 (o_0r1[3:3]);
  GND I36 (o_0r1[4:4]);
  GND I37 (o_0r1[5:5]);
  GND I38 (o_0r1[6:6]);
  GND I39 (o_0r1[7:7]);
  GND I40 (o_0r1[8:8]);
  GND I41 (o_0r1[9:9]);
  GND I42 (o_0r1[10:10]);
  GND I43 (o_0r1[11:11]);
  GND I44 (o_0r1[12:12]);
  GND I45 (o_0r1[13:13]);
  GND I46 (o_0r1[14:14]);
  GND I47 (o_0r1[15:15]);
  GND I48 (o_0r1[16:16]);
  GND I49 (o_0r1[17:17]);
  GND I50 (o_0r1[18:18]);
  GND I51 (o_0r1[19:19]);
  GND I52 (o_0r1[20:20]);
  GND I53 (o_0r1[21:21]);
  GND I54 (o_0r1[22:22]);
  GND I55 (o_0r1[23:23]);
  GND I56 (o_0r1[24:24]);
  GND I57 (o_0r1[25:25]);
  GND I58 (o_0r1[26:26]);
  GND I59 (o_0r1[27:27]);
  GND I60 (o_0r1[28:28]);
  GND I61 (o_0r1[29:29]);
  GND I62 (o_0r1[30:30]);
  GND I63 (o_0r1[31:31]);
  BUFF I64 (i_0a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0 TeakF [0,0,0] [One 0,Many [0,0,0]]
module tkf0mo0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  C3 I3 (i_0a, o_0a, o_1a, o_2a);
endmodule

// tkj0m0_0 TeakJ [Many [0,0],One 0]
module tkj0m0_0 (i_0r, i_0a, i_1r, i_1a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input reset;
  C2 I0 (o_0r, i_0r, i_1r);
  BUFF I1 (i_0a, o_0a);
  BUFF I2 (i_1a, o_0a);
endmodule

// tko0m32_1nm32b0 TeakO [
//     (1,TeakOConstant 32 0)] [One 0,One 32]
module tko0m32_1nm32b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  BUFF I6 (o_0r0[6:6], i_0r);
  BUFF I7 (o_0r0[7:7], i_0r);
  BUFF I8 (o_0r0[8:8], i_0r);
  BUFF I9 (o_0r0[9:9], i_0r);
  BUFF I10 (o_0r0[10:10], i_0r);
  BUFF I11 (o_0r0[11:11], i_0r);
  BUFF I12 (o_0r0[12:12], i_0r);
  BUFF I13 (o_0r0[13:13], i_0r);
  BUFF I14 (o_0r0[14:14], i_0r);
  BUFF I15 (o_0r0[15:15], i_0r);
  BUFF I16 (o_0r0[16:16], i_0r);
  BUFF I17 (o_0r0[17:17], i_0r);
  BUFF I18 (o_0r0[18:18], i_0r);
  BUFF I19 (o_0r0[19:19], i_0r);
  BUFF I20 (o_0r0[20:20], i_0r);
  BUFF I21 (o_0r0[21:21], i_0r);
  BUFF I22 (o_0r0[22:22], i_0r);
  BUFF I23 (o_0r0[23:23], i_0r);
  BUFF I24 (o_0r0[24:24], i_0r);
  BUFF I25 (o_0r0[25:25], i_0r);
  BUFF I26 (o_0r0[26:26], i_0r);
  BUFF I27 (o_0r0[27:27], i_0r);
  BUFF I28 (o_0r0[28:28], i_0r);
  BUFF I29 (o_0r0[29:29], i_0r);
  BUFF I30 (o_0r0[30:30], i_0r);
  BUFF I31 (o_0r0[31:31], i_0r);
  GND I32 (o_0r1[0:0]);
  GND I33 (o_0r1[1:1]);
  GND I34 (o_0r1[2:2]);
  GND I35 (o_0r1[3:3]);
  GND I36 (o_0r1[4:4]);
  GND I37 (o_0r1[5:5]);
  GND I38 (o_0r1[6:6]);
  GND I39 (o_0r1[7:7]);
  GND I40 (o_0r1[8:8]);
  GND I41 (o_0r1[9:9]);
  GND I42 (o_0r1[10:10]);
  GND I43 (o_0r1[11:11]);
  GND I44 (o_0r1[12:12]);
  GND I45 (o_0r1[13:13]);
  GND I46 (o_0r1[14:14]);
  GND I47 (o_0r1[15:15]);
  GND I48 (o_0r1[16:16]);
  GND I49 (o_0r1[17:17]);
  GND I50 (o_0r1[18:18]);
  GND I51 (o_0r1[19:19]);
  GND I52 (o_0r1[20:20]);
  GND I53 (o_0r1[21:21]);
  GND I54 (o_0r1[22:22]);
  GND I55 (o_0r1[23:23]);
  GND I56 (o_0r1[24:24]);
  GND I57 (o_0r1[25:25]);
  GND I58 (o_0r1[26:26]);
  GND I59 (o_0r1[27:27]);
  GND I60 (o_0r1[28:28]);
  GND I61 (o_0r1[29:29]);
  GND I62 (o_0r1[30:30]);
  GND I63 (o_0r1[31:31]);
  BUFF I64 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b0 TeakO [
//     (1,TeakOConstant 3 0)] [One 0,One 3]
module tko0m3_1nm3b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  GND I3 (o_0r1[0:0]);
  GND I4 (o_0r1[1:1]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko32m32_1nm32b0_2subt1o0w32bi0w32b TeakO [
//     (1,TeakOConstant 32 0),
//     (2,TeakOp TeakOpSub [(1,0+:32),(0,0+:32)])] [One 32,One 32]
module tko32m32_1nm32b0_2subt1o0w32bi0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [31:0] gocomp_0;
  wire [10:0] simp341_0;
  wire [3:0] simp342_0;
  wire [1:0] simp343_0;
  wire [31:0] termf_1;
  wire [31:0] termt_1;
  wire [31:0] cf2__0;
  wire [31:0] ct2__0;
  wire [3:0] ha2__0;
  wire [7:0] fa2_1min_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [7:0] fa2_2min_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  wire [7:0] fa2_3min_0;
  wire [1:0] simp861_0;
  wire [1:0] simp871_0;
  wire [7:0] fa2_4min_0;
  wire [1:0] simp991_0;
  wire [1:0] simp1001_0;
  wire [7:0] fa2_5min_0;
  wire [1:0] simp1121_0;
  wire [1:0] simp1131_0;
  wire [7:0] fa2_6min_0;
  wire [1:0] simp1251_0;
  wire [1:0] simp1261_0;
  wire [7:0] fa2_7min_0;
  wire [1:0] simp1381_0;
  wire [1:0] simp1391_0;
  wire [7:0] fa2_8min_0;
  wire [1:0] simp1511_0;
  wire [1:0] simp1521_0;
  wire [7:0] fa2_9min_0;
  wire [1:0] simp1641_0;
  wire [1:0] simp1651_0;
  wire [7:0] fa2_10min_0;
  wire [1:0] simp1771_0;
  wire [1:0] simp1781_0;
  wire [7:0] fa2_11min_0;
  wire [1:0] simp1901_0;
  wire [1:0] simp1911_0;
  wire [7:0] fa2_12min_0;
  wire [1:0] simp2031_0;
  wire [1:0] simp2041_0;
  wire [7:0] fa2_13min_0;
  wire [1:0] simp2161_0;
  wire [1:0] simp2171_0;
  wire [7:0] fa2_14min_0;
  wire [1:0] simp2291_0;
  wire [1:0] simp2301_0;
  wire [7:0] fa2_15min_0;
  wire [1:0] simp2421_0;
  wire [1:0] simp2431_0;
  wire [7:0] fa2_16min_0;
  wire [1:0] simp2551_0;
  wire [1:0] simp2561_0;
  wire [7:0] fa2_17min_0;
  wire [1:0] simp2681_0;
  wire [1:0] simp2691_0;
  wire [7:0] fa2_18min_0;
  wire [1:0] simp2811_0;
  wire [1:0] simp2821_0;
  wire [7:0] fa2_19min_0;
  wire [1:0] simp2941_0;
  wire [1:0] simp2951_0;
  wire [7:0] fa2_20min_0;
  wire [1:0] simp3071_0;
  wire [1:0] simp3081_0;
  wire [7:0] fa2_21min_0;
  wire [1:0] simp3201_0;
  wire [1:0] simp3211_0;
  wire [7:0] fa2_22min_0;
  wire [1:0] simp3331_0;
  wire [1:0] simp3341_0;
  wire [7:0] fa2_23min_0;
  wire [1:0] simp3461_0;
  wire [1:0] simp3471_0;
  wire [7:0] fa2_24min_0;
  wire [1:0] simp3591_0;
  wire [1:0] simp3601_0;
  wire [7:0] fa2_25min_0;
  wire [1:0] simp3721_0;
  wire [1:0] simp3731_0;
  wire [7:0] fa2_26min_0;
  wire [1:0] simp3851_0;
  wire [1:0] simp3861_0;
  wire [7:0] fa2_27min_0;
  wire [1:0] simp3981_0;
  wire [1:0] simp3991_0;
  wire [7:0] fa2_28min_0;
  wire [1:0] simp4111_0;
  wire [1:0] simp4121_0;
  wire [7:0] fa2_29min_0;
  wire [1:0] simp4241_0;
  wire [1:0] simp4251_0;
  wire [7:0] fa2_30min_0;
  wire [1:0] simp4371_0;
  wire [1:0] simp4381_0;
  wire [7:0] fa2_31min_0;
  wire [1:0] simp4501_0;
  wire [1:0] simp4511_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I32 (simp341_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I33 (simp341_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I34 (simp341_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I35 (simp341_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I36 (simp341_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I37 (simp341_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I38 (simp341_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I39 (simp341_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I40 (simp341_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I41 (simp341_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C2 I42 (simp341_0[10:10], gocomp_0[30:30], gocomp_0[31:31]);
  C3 I43 (simp342_0[0:0], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  C3 I44 (simp342_0[1:1], simp341_0[3:3], simp341_0[4:4], simp341_0[5:5]);
  C3 I45 (simp342_0[2:2], simp341_0[6:6], simp341_0[7:7], simp341_0[8:8]);
  C2 I46 (simp342_0[3:3], simp341_0[9:9], simp341_0[10:10]);
  C3 I47 (simp343_0[0:0], simp342_0[0:0], simp342_0[1:1], simp342_0[2:2]);
  BUFF I48 (simp343_0[1:1], simp342_0[3:3]);
  C2 I49 (go_0, simp343_0[0:0], simp343_0[1:1]);
  BUFF I50 (termf_1[0:0], go_0);
  BUFF I51 (termf_1[1:1], go_0);
  BUFF I52 (termf_1[2:2], go_0);
  BUFF I53 (termf_1[3:3], go_0);
  BUFF I54 (termf_1[4:4], go_0);
  BUFF I55 (termf_1[5:5], go_0);
  BUFF I56 (termf_1[6:6], go_0);
  BUFF I57 (termf_1[7:7], go_0);
  BUFF I58 (termf_1[8:8], go_0);
  BUFF I59 (termf_1[9:9], go_0);
  BUFF I60 (termf_1[10:10], go_0);
  BUFF I61 (termf_1[11:11], go_0);
  BUFF I62 (termf_1[12:12], go_0);
  BUFF I63 (termf_1[13:13], go_0);
  BUFF I64 (termf_1[14:14], go_0);
  BUFF I65 (termf_1[15:15], go_0);
  BUFF I66 (termf_1[16:16], go_0);
  BUFF I67 (termf_1[17:17], go_0);
  BUFF I68 (termf_1[18:18], go_0);
  BUFF I69 (termf_1[19:19], go_0);
  BUFF I70 (termf_1[20:20], go_0);
  BUFF I71 (termf_1[21:21], go_0);
  BUFF I72 (termf_1[22:22], go_0);
  BUFF I73 (termf_1[23:23], go_0);
  BUFF I74 (termf_1[24:24], go_0);
  BUFF I75 (termf_1[25:25], go_0);
  BUFF I76 (termf_1[26:26], go_0);
  BUFF I77 (termf_1[27:27], go_0);
  BUFF I78 (termf_1[28:28], go_0);
  BUFF I79 (termf_1[29:29], go_0);
  BUFF I80 (termf_1[30:30], go_0);
  BUFF I81 (termf_1[31:31], go_0);
  GND I82 (termt_1[0:0]);
  GND I83 (termt_1[1:1]);
  GND I84 (termt_1[2:2]);
  GND I85 (termt_1[3:3]);
  GND I86 (termt_1[4:4]);
  GND I87 (termt_1[5:5]);
  GND I88 (termt_1[6:6]);
  GND I89 (termt_1[7:7]);
  GND I90 (termt_1[8:8]);
  GND I91 (termt_1[9:9]);
  GND I92 (termt_1[10:10]);
  GND I93 (termt_1[11:11]);
  GND I94 (termt_1[12:12]);
  GND I95 (termt_1[13:13]);
  GND I96 (termt_1[14:14]);
  GND I97 (termt_1[15:15]);
  GND I98 (termt_1[16:16]);
  GND I99 (termt_1[17:17]);
  GND I100 (termt_1[18:18]);
  GND I101 (termt_1[19:19]);
  GND I102 (termt_1[20:20]);
  GND I103 (termt_1[21:21]);
  GND I104 (termt_1[22:22]);
  GND I105 (termt_1[23:23]);
  GND I106 (termt_1[24:24]);
  GND I107 (termt_1[25:25]);
  GND I108 (termt_1[26:26]);
  GND I109 (termt_1[27:27]);
  GND I110 (termt_1[28:28]);
  GND I111 (termt_1[29:29]);
  GND I112 (termt_1[30:30]);
  GND I113 (termt_1[31:31]);
  C2 I114 (ha2__0[0:0], i_0r1[0:0], termf_1[0:0]);
  C2 I115 (ha2__0[1:1], i_0r1[0:0], termt_1[0:0]);
  C2 I116 (ha2__0[2:2], i_0r0[0:0], termf_1[0:0]);
  C2 I117 (ha2__0[3:3], i_0r0[0:0], termt_1[0:0]);
  BUFF I118 (cf2__0[0:0], ha2__0[0:0]);
  OR3 I119 (ct2__0[0:0], ha2__0[1:1], ha2__0[2:2], ha2__0[3:3]);
  OR2 I120 (o_0r0[0:0], ha2__0[1:1], ha2__0[2:2]);
  OR2 I121 (o_0r1[0:0], ha2__0[0:0], ha2__0[3:3]);
  C3 I122 (fa2_1min_0[0:0], cf2__0[0:0], i_0r1[1:1], termf_1[1:1]);
  C3 I123 (fa2_1min_0[1:1], cf2__0[0:0], i_0r1[1:1], termt_1[1:1]);
  C3 I124 (fa2_1min_0[2:2], cf2__0[0:0], i_0r0[1:1], termf_1[1:1]);
  C3 I125 (fa2_1min_0[3:3], cf2__0[0:0], i_0r0[1:1], termt_1[1:1]);
  C3 I126 (fa2_1min_0[4:4], ct2__0[0:0], i_0r1[1:1], termf_1[1:1]);
  C3 I127 (fa2_1min_0[5:5], ct2__0[0:0], i_0r1[1:1], termt_1[1:1]);
  C3 I128 (fa2_1min_0[6:6], ct2__0[0:0], i_0r0[1:1], termf_1[1:1]);
  C3 I129 (fa2_1min_0[7:7], ct2__0[0:0], i_0r0[1:1], termt_1[1:1]);
  NOR3 I130 (simp601_0[0:0], fa2_1min_0[0:0], fa2_1min_0[3:3], fa2_1min_0[5:5]);
  INV I131 (simp601_0[1:1], fa2_1min_0[6:6]);
  NAND2 I132 (o_0r0[1:1], simp601_0[0:0], simp601_0[1:1]);
  NOR3 I133 (simp611_0[0:0], fa2_1min_0[1:1], fa2_1min_0[2:2], fa2_1min_0[4:4]);
  INV I134 (simp611_0[1:1], fa2_1min_0[7:7]);
  NAND2 I135 (o_0r1[1:1], simp611_0[0:0], simp611_0[1:1]);
  AO222 I136 (ct2__0[1:1], termt_1[1:1], i_0r0[1:1], termt_1[1:1], ct2__0[0:0], i_0r0[1:1], ct2__0[0:0]);
  AO222 I137 (cf2__0[1:1], termf_1[1:1], i_0r1[1:1], termf_1[1:1], cf2__0[0:0], i_0r1[1:1], cf2__0[0:0]);
  C3 I138 (fa2_2min_0[0:0], cf2__0[1:1], i_0r1[2:2], termf_1[2:2]);
  C3 I139 (fa2_2min_0[1:1], cf2__0[1:1], i_0r1[2:2], termt_1[2:2]);
  C3 I140 (fa2_2min_0[2:2], cf2__0[1:1], i_0r0[2:2], termf_1[2:2]);
  C3 I141 (fa2_2min_0[3:3], cf2__0[1:1], i_0r0[2:2], termt_1[2:2]);
  C3 I142 (fa2_2min_0[4:4], ct2__0[1:1], i_0r1[2:2], termf_1[2:2]);
  C3 I143 (fa2_2min_0[5:5], ct2__0[1:1], i_0r1[2:2], termt_1[2:2]);
  C3 I144 (fa2_2min_0[6:6], ct2__0[1:1], i_0r0[2:2], termf_1[2:2]);
  C3 I145 (fa2_2min_0[7:7], ct2__0[1:1], i_0r0[2:2], termt_1[2:2]);
  NOR3 I146 (simp731_0[0:0], fa2_2min_0[0:0], fa2_2min_0[3:3], fa2_2min_0[5:5]);
  INV I147 (simp731_0[1:1], fa2_2min_0[6:6]);
  NAND2 I148 (o_0r0[2:2], simp731_0[0:0], simp731_0[1:1]);
  NOR3 I149 (simp741_0[0:0], fa2_2min_0[1:1], fa2_2min_0[2:2], fa2_2min_0[4:4]);
  INV I150 (simp741_0[1:1], fa2_2min_0[7:7]);
  NAND2 I151 (o_0r1[2:2], simp741_0[0:0], simp741_0[1:1]);
  AO222 I152 (ct2__0[2:2], termt_1[2:2], i_0r0[2:2], termt_1[2:2], ct2__0[1:1], i_0r0[2:2], ct2__0[1:1]);
  AO222 I153 (cf2__0[2:2], termf_1[2:2], i_0r1[2:2], termf_1[2:2], cf2__0[1:1], i_0r1[2:2], cf2__0[1:1]);
  C3 I154 (fa2_3min_0[0:0], cf2__0[2:2], i_0r1[3:3], termf_1[3:3]);
  C3 I155 (fa2_3min_0[1:1], cf2__0[2:2], i_0r1[3:3], termt_1[3:3]);
  C3 I156 (fa2_3min_0[2:2], cf2__0[2:2], i_0r0[3:3], termf_1[3:3]);
  C3 I157 (fa2_3min_0[3:3], cf2__0[2:2], i_0r0[3:3], termt_1[3:3]);
  C3 I158 (fa2_3min_0[4:4], ct2__0[2:2], i_0r1[3:3], termf_1[3:3]);
  C3 I159 (fa2_3min_0[5:5], ct2__0[2:2], i_0r1[3:3], termt_1[3:3]);
  C3 I160 (fa2_3min_0[6:6], ct2__0[2:2], i_0r0[3:3], termf_1[3:3]);
  C3 I161 (fa2_3min_0[7:7], ct2__0[2:2], i_0r0[3:3], termt_1[3:3]);
  NOR3 I162 (simp861_0[0:0], fa2_3min_0[0:0], fa2_3min_0[3:3], fa2_3min_0[5:5]);
  INV I163 (simp861_0[1:1], fa2_3min_0[6:6]);
  NAND2 I164 (o_0r0[3:3], simp861_0[0:0], simp861_0[1:1]);
  NOR3 I165 (simp871_0[0:0], fa2_3min_0[1:1], fa2_3min_0[2:2], fa2_3min_0[4:4]);
  INV I166 (simp871_0[1:1], fa2_3min_0[7:7]);
  NAND2 I167 (o_0r1[3:3], simp871_0[0:0], simp871_0[1:1]);
  AO222 I168 (ct2__0[3:3], termt_1[3:3], i_0r0[3:3], termt_1[3:3], ct2__0[2:2], i_0r0[3:3], ct2__0[2:2]);
  AO222 I169 (cf2__0[3:3], termf_1[3:3], i_0r1[3:3], termf_1[3:3], cf2__0[2:2], i_0r1[3:3], cf2__0[2:2]);
  C3 I170 (fa2_4min_0[0:0], cf2__0[3:3], i_0r1[4:4], termf_1[4:4]);
  C3 I171 (fa2_4min_0[1:1], cf2__0[3:3], i_0r1[4:4], termt_1[4:4]);
  C3 I172 (fa2_4min_0[2:2], cf2__0[3:3], i_0r0[4:4], termf_1[4:4]);
  C3 I173 (fa2_4min_0[3:3], cf2__0[3:3], i_0r0[4:4], termt_1[4:4]);
  C3 I174 (fa2_4min_0[4:4], ct2__0[3:3], i_0r1[4:4], termf_1[4:4]);
  C3 I175 (fa2_4min_0[5:5], ct2__0[3:3], i_0r1[4:4], termt_1[4:4]);
  C3 I176 (fa2_4min_0[6:6], ct2__0[3:3], i_0r0[4:4], termf_1[4:4]);
  C3 I177 (fa2_4min_0[7:7], ct2__0[3:3], i_0r0[4:4], termt_1[4:4]);
  NOR3 I178 (simp991_0[0:0], fa2_4min_0[0:0], fa2_4min_0[3:3], fa2_4min_0[5:5]);
  INV I179 (simp991_0[1:1], fa2_4min_0[6:6]);
  NAND2 I180 (o_0r0[4:4], simp991_0[0:0], simp991_0[1:1]);
  NOR3 I181 (simp1001_0[0:0], fa2_4min_0[1:1], fa2_4min_0[2:2], fa2_4min_0[4:4]);
  INV I182 (simp1001_0[1:1], fa2_4min_0[7:7]);
  NAND2 I183 (o_0r1[4:4], simp1001_0[0:0], simp1001_0[1:1]);
  AO222 I184 (ct2__0[4:4], termt_1[4:4], i_0r0[4:4], termt_1[4:4], ct2__0[3:3], i_0r0[4:4], ct2__0[3:3]);
  AO222 I185 (cf2__0[4:4], termf_1[4:4], i_0r1[4:4], termf_1[4:4], cf2__0[3:3], i_0r1[4:4], cf2__0[3:3]);
  C3 I186 (fa2_5min_0[0:0], cf2__0[4:4], i_0r1[5:5], termf_1[5:5]);
  C3 I187 (fa2_5min_0[1:1], cf2__0[4:4], i_0r1[5:5], termt_1[5:5]);
  C3 I188 (fa2_5min_0[2:2], cf2__0[4:4], i_0r0[5:5], termf_1[5:5]);
  C3 I189 (fa2_5min_0[3:3], cf2__0[4:4], i_0r0[5:5], termt_1[5:5]);
  C3 I190 (fa2_5min_0[4:4], ct2__0[4:4], i_0r1[5:5], termf_1[5:5]);
  C3 I191 (fa2_5min_0[5:5], ct2__0[4:4], i_0r1[5:5], termt_1[5:5]);
  C3 I192 (fa2_5min_0[6:6], ct2__0[4:4], i_0r0[5:5], termf_1[5:5]);
  C3 I193 (fa2_5min_0[7:7], ct2__0[4:4], i_0r0[5:5], termt_1[5:5]);
  NOR3 I194 (simp1121_0[0:0], fa2_5min_0[0:0], fa2_5min_0[3:3], fa2_5min_0[5:5]);
  INV I195 (simp1121_0[1:1], fa2_5min_0[6:6]);
  NAND2 I196 (o_0r0[5:5], simp1121_0[0:0], simp1121_0[1:1]);
  NOR3 I197 (simp1131_0[0:0], fa2_5min_0[1:1], fa2_5min_0[2:2], fa2_5min_0[4:4]);
  INV I198 (simp1131_0[1:1], fa2_5min_0[7:7]);
  NAND2 I199 (o_0r1[5:5], simp1131_0[0:0], simp1131_0[1:1]);
  AO222 I200 (ct2__0[5:5], termt_1[5:5], i_0r0[5:5], termt_1[5:5], ct2__0[4:4], i_0r0[5:5], ct2__0[4:4]);
  AO222 I201 (cf2__0[5:5], termf_1[5:5], i_0r1[5:5], termf_1[5:5], cf2__0[4:4], i_0r1[5:5], cf2__0[4:4]);
  C3 I202 (fa2_6min_0[0:0], cf2__0[5:5], i_0r1[6:6], termf_1[6:6]);
  C3 I203 (fa2_6min_0[1:1], cf2__0[5:5], i_0r1[6:6], termt_1[6:6]);
  C3 I204 (fa2_6min_0[2:2], cf2__0[5:5], i_0r0[6:6], termf_1[6:6]);
  C3 I205 (fa2_6min_0[3:3], cf2__0[5:5], i_0r0[6:6], termt_1[6:6]);
  C3 I206 (fa2_6min_0[4:4], ct2__0[5:5], i_0r1[6:6], termf_1[6:6]);
  C3 I207 (fa2_6min_0[5:5], ct2__0[5:5], i_0r1[6:6], termt_1[6:6]);
  C3 I208 (fa2_6min_0[6:6], ct2__0[5:5], i_0r0[6:6], termf_1[6:6]);
  C3 I209 (fa2_6min_0[7:7], ct2__0[5:5], i_0r0[6:6], termt_1[6:6]);
  NOR3 I210 (simp1251_0[0:0], fa2_6min_0[0:0], fa2_6min_0[3:3], fa2_6min_0[5:5]);
  INV I211 (simp1251_0[1:1], fa2_6min_0[6:6]);
  NAND2 I212 (o_0r0[6:6], simp1251_0[0:0], simp1251_0[1:1]);
  NOR3 I213 (simp1261_0[0:0], fa2_6min_0[1:1], fa2_6min_0[2:2], fa2_6min_0[4:4]);
  INV I214 (simp1261_0[1:1], fa2_6min_0[7:7]);
  NAND2 I215 (o_0r1[6:6], simp1261_0[0:0], simp1261_0[1:1]);
  AO222 I216 (ct2__0[6:6], termt_1[6:6], i_0r0[6:6], termt_1[6:6], ct2__0[5:5], i_0r0[6:6], ct2__0[5:5]);
  AO222 I217 (cf2__0[6:6], termf_1[6:6], i_0r1[6:6], termf_1[6:6], cf2__0[5:5], i_0r1[6:6], cf2__0[5:5]);
  C3 I218 (fa2_7min_0[0:0], cf2__0[6:6], i_0r1[7:7], termf_1[7:7]);
  C3 I219 (fa2_7min_0[1:1], cf2__0[6:6], i_0r1[7:7], termt_1[7:7]);
  C3 I220 (fa2_7min_0[2:2], cf2__0[6:6], i_0r0[7:7], termf_1[7:7]);
  C3 I221 (fa2_7min_0[3:3], cf2__0[6:6], i_0r0[7:7], termt_1[7:7]);
  C3 I222 (fa2_7min_0[4:4], ct2__0[6:6], i_0r1[7:7], termf_1[7:7]);
  C3 I223 (fa2_7min_0[5:5], ct2__0[6:6], i_0r1[7:7], termt_1[7:7]);
  C3 I224 (fa2_7min_0[6:6], ct2__0[6:6], i_0r0[7:7], termf_1[7:7]);
  C3 I225 (fa2_7min_0[7:7], ct2__0[6:6], i_0r0[7:7], termt_1[7:7]);
  NOR3 I226 (simp1381_0[0:0], fa2_7min_0[0:0], fa2_7min_0[3:3], fa2_7min_0[5:5]);
  INV I227 (simp1381_0[1:1], fa2_7min_0[6:6]);
  NAND2 I228 (o_0r0[7:7], simp1381_0[0:0], simp1381_0[1:1]);
  NOR3 I229 (simp1391_0[0:0], fa2_7min_0[1:1], fa2_7min_0[2:2], fa2_7min_0[4:4]);
  INV I230 (simp1391_0[1:1], fa2_7min_0[7:7]);
  NAND2 I231 (o_0r1[7:7], simp1391_0[0:0], simp1391_0[1:1]);
  AO222 I232 (ct2__0[7:7], termt_1[7:7], i_0r0[7:7], termt_1[7:7], ct2__0[6:6], i_0r0[7:7], ct2__0[6:6]);
  AO222 I233 (cf2__0[7:7], termf_1[7:7], i_0r1[7:7], termf_1[7:7], cf2__0[6:6], i_0r1[7:7], cf2__0[6:6]);
  C3 I234 (fa2_8min_0[0:0], cf2__0[7:7], i_0r1[8:8], termf_1[8:8]);
  C3 I235 (fa2_8min_0[1:1], cf2__0[7:7], i_0r1[8:8], termt_1[8:8]);
  C3 I236 (fa2_8min_0[2:2], cf2__0[7:7], i_0r0[8:8], termf_1[8:8]);
  C3 I237 (fa2_8min_0[3:3], cf2__0[7:7], i_0r0[8:8], termt_1[8:8]);
  C3 I238 (fa2_8min_0[4:4], ct2__0[7:7], i_0r1[8:8], termf_1[8:8]);
  C3 I239 (fa2_8min_0[5:5], ct2__0[7:7], i_0r1[8:8], termt_1[8:8]);
  C3 I240 (fa2_8min_0[6:6], ct2__0[7:7], i_0r0[8:8], termf_1[8:8]);
  C3 I241 (fa2_8min_0[7:7], ct2__0[7:7], i_0r0[8:8], termt_1[8:8]);
  NOR3 I242 (simp1511_0[0:0], fa2_8min_0[0:0], fa2_8min_0[3:3], fa2_8min_0[5:5]);
  INV I243 (simp1511_0[1:1], fa2_8min_0[6:6]);
  NAND2 I244 (o_0r0[8:8], simp1511_0[0:0], simp1511_0[1:1]);
  NOR3 I245 (simp1521_0[0:0], fa2_8min_0[1:1], fa2_8min_0[2:2], fa2_8min_0[4:4]);
  INV I246 (simp1521_0[1:1], fa2_8min_0[7:7]);
  NAND2 I247 (o_0r1[8:8], simp1521_0[0:0], simp1521_0[1:1]);
  AO222 I248 (ct2__0[8:8], termt_1[8:8], i_0r0[8:8], termt_1[8:8], ct2__0[7:7], i_0r0[8:8], ct2__0[7:7]);
  AO222 I249 (cf2__0[8:8], termf_1[8:8], i_0r1[8:8], termf_1[8:8], cf2__0[7:7], i_0r1[8:8], cf2__0[7:7]);
  C3 I250 (fa2_9min_0[0:0], cf2__0[8:8], i_0r1[9:9], termf_1[9:9]);
  C3 I251 (fa2_9min_0[1:1], cf2__0[8:8], i_0r1[9:9], termt_1[9:9]);
  C3 I252 (fa2_9min_0[2:2], cf2__0[8:8], i_0r0[9:9], termf_1[9:9]);
  C3 I253 (fa2_9min_0[3:3], cf2__0[8:8], i_0r0[9:9], termt_1[9:9]);
  C3 I254 (fa2_9min_0[4:4], ct2__0[8:8], i_0r1[9:9], termf_1[9:9]);
  C3 I255 (fa2_9min_0[5:5], ct2__0[8:8], i_0r1[9:9], termt_1[9:9]);
  C3 I256 (fa2_9min_0[6:6], ct2__0[8:8], i_0r0[9:9], termf_1[9:9]);
  C3 I257 (fa2_9min_0[7:7], ct2__0[8:8], i_0r0[9:9], termt_1[9:9]);
  NOR3 I258 (simp1641_0[0:0], fa2_9min_0[0:0], fa2_9min_0[3:3], fa2_9min_0[5:5]);
  INV I259 (simp1641_0[1:1], fa2_9min_0[6:6]);
  NAND2 I260 (o_0r0[9:9], simp1641_0[0:0], simp1641_0[1:1]);
  NOR3 I261 (simp1651_0[0:0], fa2_9min_0[1:1], fa2_9min_0[2:2], fa2_9min_0[4:4]);
  INV I262 (simp1651_0[1:1], fa2_9min_0[7:7]);
  NAND2 I263 (o_0r1[9:9], simp1651_0[0:0], simp1651_0[1:1]);
  AO222 I264 (ct2__0[9:9], termt_1[9:9], i_0r0[9:9], termt_1[9:9], ct2__0[8:8], i_0r0[9:9], ct2__0[8:8]);
  AO222 I265 (cf2__0[9:9], termf_1[9:9], i_0r1[9:9], termf_1[9:9], cf2__0[8:8], i_0r1[9:9], cf2__0[8:8]);
  C3 I266 (fa2_10min_0[0:0], cf2__0[9:9], i_0r1[10:10], termf_1[10:10]);
  C3 I267 (fa2_10min_0[1:1], cf2__0[9:9], i_0r1[10:10], termt_1[10:10]);
  C3 I268 (fa2_10min_0[2:2], cf2__0[9:9], i_0r0[10:10], termf_1[10:10]);
  C3 I269 (fa2_10min_0[3:3], cf2__0[9:9], i_0r0[10:10], termt_1[10:10]);
  C3 I270 (fa2_10min_0[4:4], ct2__0[9:9], i_0r1[10:10], termf_1[10:10]);
  C3 I271 (fa2_10min_0[5:5], ct2__0[9:9], i_0r1[10:10], termt_1[10:10]);
  C3 I272 (fa2_10min_0[6:6], ct2__0[9:9], i_0r0[10:10], termf_1[10:10]);
  C3 I273 (fa2_10min_0[7:7], ct2__0[9:9], i_0r0[10:10], termt_1[10:10]);
  NOR3 I274 (simp1771_0[0:0], fa2_10min_0[0:0], fa2_10min_0[3:3], fa2_10min_0[5:5]);
  INV I275 (simp1771_0[1:1], fa2_10min_0[6:6]);
  NAND2 I276 (o_0r0[10:10], simp1771_0[0:0], simp1771_0[1:1]);
  NOR3 I277 (simp1781_0[0:0], fa2_10min_0[1:1], fa2_10min_0[2:2], fa2_10min_0[4:4]);
  INV I278 (simp1781_0[1:1], fa2_10min_0[7:7]);
  NAND2 I279 (o_0r1[10:10], simp1781_0[0:0], simp1781_0[1:1]);
  AO222 I280 (ct2__0[10:10], termt_1[10:10], i_0r0[10:10], termt_1[10:10], ct2__0[9:9], i_0r0[10:10], ct2__0[9:9]);
  AO222 I281 (cf2__0[10:10], termf_1[10:10], i_0r1[10:10], termf_1[10:10], cf2__0[9:9], i_0r1[10:10], cf2__0[9:9]);
  C3 I282 (fa2_11min_0[0:0], cf2__0[10:10], i_0r1[11:11], termf_1[11:11]);
  C3 I283 (fa2_11min_0[1:1], cf2__0[10:10], i_0r1[11:11], termt_1[11:11]);
  C3 I284 (fa2_11min_0[2:2], cf2__0[10:10], i_0r0[11:11], termf_1[11:11]);
  C3 I285 (fa2_11min_0[3:3], cf2__0[10:10], i_0r0[11:11], termt_1[11:11]);
  C3 I286 (fa2_11min_0[4:4], ct2__0[10:10], i_0r1[11:11], termf_1[11:11]);
  C3 I287 (fa2_11min_0[5:5], ct2__0[10:10], i_0r1[11:11], termt_1[11:11]);
  C3 I288 (fa2_11min_0[6:6], ct2__0[10:10], i_0r0[11:11], termf_1[11:11]);
  C3 I289 (fa2_11min_0[7:7], ct2__0[10:10], i_0r0[11:11], termt_1[11:11]);
  NOR3 I290 (simp1901_0[0:0], fa2_11min_0[0:0], fa2_11min_0[3:3], fa2_11min_0[5:5]);
  INV I291 (simp1901_0[1:1], fa2_11min_0[6:6]);
  NAND2 I292 (o_0r0[11:11], simp1901_0[0:0], simp1901_0[1:1]);
  NOR3 I293 (simp1911_0[0:0], fa2_11min_0[1:1], fa2_11min_0[2:2], fa2_11min_0[4:4]);
  INV I294 (simp1911_0[1:1], fa2_11min_0[7:7]);
  NAND2 I295 (o_0r1[11:11], simp1911_0[0:0], simp1911_0[1:1]);
  AO222 I296 (ct2__0[11:11], termt_1[11:11], i_0r0[11:11], termt_1[11:11], ct2__0[10:10], i_0r0[11:11], ct2__0[10:10]);
  AO222 I297 (cf2__0[11:11], termf_1[11:11], i_0r1[11:11], termf_1[11:11], cf2__0[10:10], i_0r1[11:11], cf2__0[10:10]);
  C3 I298 (fa2_12min_0[0:0], cf2__0[11:11], i_0r1[12:12], termf_1[12:12]);
  C3 I299 (fa2_12min_0[1:1], cf2__0[11:11], i_0r1[12:12], termt_1[12:12]);
  C3 I300 (fa2_12min_0[2:2], cf2__0[11:11], i_0r0[12:12], termf_1[12:12]);
  C3 I301 (fa2_12min_0[3:3], cf2__0[11:11], i_0r0[12:12], termt_1[12:12]);
  C3 I302 (fa2_12min_0[4:4], ct2__0[11:11], i_0r1[12:12], termf_1[12:12]);
  C3 I303 (fa2_12min_0[5:5], ct2__0[11:11], i_0r1[12:12], termt_1[12:12]);
  C3 I304 (fa2_12min_0[6:6], ct2__0[11:11], i_0r0[12:12], termf_1[12:12]);
  C3 I305 (fa2_12min_0[7:7], ct2__0[11:11], i_0r0[12:12], termt_1[12:12]);
  NOR3 I306 (simp2031_0[0:0], fa2_12min_0[0:0], fa2_12min_0[3:3], fa2_12min_0[5:5]);
  INV I307 (simp2031_0[1:1], fa2_12min_0[6:6]);
  NAND2 I308 (o_0r0[12:12], simp2031_0[0:0], simp2031_0[1:1]);
  NOR3 I309 (simp2041_0[0:0], fa2_12min_0[1:1], fa2_12min_0[2:2], fa2_12min_0[4:4]);
  INV I310 (simp2041_0[1:1], fa2_12min_0[7:7]);
  NAND2 I311 (o_0r1[12:12], simp2041_0[0:0], simp2041_0[1:1]);
  AO222 I312 (ct2__0[12:12], termt_1[12:12], i_0r0[12:12], termt_1[12:12], ct2__0[11:11], i_0r0[12:12], ct2__0[11:11]);
  AO222 I313 (cf2__0[12:12], termf_1[12:12], i_0r1[12:12], termf_1[12:12], cf2__0[11:11], i_0r1[12:12], cf2__0[11:11]);
  C3 I314 (fa2_13min_0[0:0], cf2__0[12:12], i_0r1[13:13], termf_1[13:13]);
  C3 I315 (fa2_13min_0[1:1], cf2__0[12:12], i_0r1[13:13], termt_1[13:13]);
  C3 I316 (fa2_13min_0[2:2], cf2__0[12:12], i_0r0[13:13], termf_1[13:13]);
  C3 I317 (fa2_13min_0[3:3], cf2__0[12:12], i_0r0[13:13], termt_1[13:13]);
  C3 I318 (fa2_13min_0[4:4], ct2__0[12:12], i_0r1[13:13], termf_1[13:13]);
  C3 I319 (fa2_13min_0[5:5], ct2__0[12:12], i_0r1[13:13], termt_1[13:13]);
  C3 I320 (fa2_13min_0[6:6], ct2__0[12:12], i_0r0[13:13], termf_1[13:13]);
  C3 I321 (fa2_13min_0[7:7], ct2__0[12:12], i_0r0[13:13], termt_1[13:13]);
  NOR3 I322 (simp2161_0[0:0], fa2_13min_0[0:0], fa2_13min_0[3:3], fa2_13min_0[5:5]);
  INV I323 (simp2161_0[1:1], fa2_13min_0[6:6]);
  NAND2 I324 (o_0r0[13:13], simp2161_0[0:0], simp2161_0[1:1]);
  NOR3 I325 (simp2171_0[0:0], fa2_13min_0[1:1], fa2_13min_0[2:2], fa2_13min_0[4:4]);
  INV I326 (simp2171_0[1:1], fa2_13min_0[7:7]);
  NAND2 I327 (o_0r1[13:13], simp2171_0[0:0], simp2171_0[1:1]);
  AO222 I328 (ct2__0[13:13], termt_1[13:13], i_0r0[13:13], termt_1[13:13], ct2__0[12:12], i_0r0[13:13], ct2__0[12:12]);
  AO222 I329 (cf2__0[13:13], termf_1[13:13], i_0r1[13:13], termf_1[13:13], cf2__0[12:12], i_0r1[13:13], cf2__0[12:12]);
  C3 I330 (fa2_14min_0[0:0], cf2__0[13:13], i_0r1[14:14], termf_1[14:14]);
  C3 I331 (fa2_14min_0[1:1], cf2__0[13:13], i_0r1[14:14], termt_1[14:14]);
  C3 I332 (fa2_14min_0[2:2], cf2__0[13:13], i_0r0[14:14], termf_1[14:14]);
  C3 I333 (fa2_14min_0[3:3], cf2__0[13:13], i_0r0[14:14], termt_1[14:14]);
  C3 I334 (fa2_14min_0[4:4], ct2__0[13:13], i_0r1[14:14], termf_1[14:14]);
  C3 I335 (fa2_14min_0[5:5], ct2__0[13:13], i_0r1[14:14], termt_1[14:14]);
  C3 I336 (fa2_14min_0[6:6], ct2__0[13:13], i_0r0[14:14], termf_1[14:14]);
  C3 I337 (fa2_14min_0[7:7], ct2__0[13:13], i_0r0[14:14], termt_1[14:14]);
  NOR3 I338 (simp2291_0[0:0], fa2_14min_0[0:0], fa2_14min_0[3:3], fa2_14min_0[5:5]);
  INV I339 (simp2291_0[1:1], fa2_14min_0[6:6]);
  NAND2 I340 (o_0r0[14:14], simp2291_0[0:0], simp2291_0[1:1]);
  NOR3 I341 (simp2301_0[0:0], fa2_14min_0[1:1], fa2_14min_0[2:2], fa2_14min_0[4:4]);
  INV I342 (simp2301_0[1:1], fa2_14min_0[7:7]);
  NAND2 I343 (o_0r1[14:14], simp2301_0[0:0], simp2301_0[1:1]);
  AO222 I344 (ct2__0[14:14], termt_1[14:14], i_0r0[14:14], termt_1[14:14], ct2__0[13:13], i_0r0[14:14], ct2__0[13:13]);
  AO222 I345 (cf2__0[14:14], termf_1[14:14], i_0r1[14:14], termf_1[14:14], cf2__0[13:13], i_0r1[14:14], cf2__0[13:13]);
  C3 I346 (fa2_15min_0[0:0], cf2__0[14:14], i_0r1[15:15], termf_1[15:15]);
  C3 I347 (fa2_15min_0[1:1], cf2__0[14:14], i_0r1[15:15], termt_1[15:15]);
  C3 I348 (fa2_15min_0[2:2], cf2__0[14:14], i_0r0[15:15], termf_1[15:15]);
  C3 I349 (fa2_15min_0[3:3], cf2__0[14:14], i_0r0[15:15], termt_1[15:15]);
  C3 I350 (fa2_15min_0[4:4], ct2__0[14:14], i_0r1[15:15], termf_1[15:15]);
  C3 I351 (fa2_15min_0[5:5], ct2__0[14:14], i_0r1[15:15], termt_1[15:15]);
  C3 I352 (fa2_15min_0[6:6], ct2__0[14:14], i_0r0[15:15], termf_1[15:15]);
  C3 I353 (fa2_15min_0[7:7], ct2__0[14:14], i_0r0[15:15], termt_1[15:15]);
  NOR3 I354 (simp2421_0[0:0], fa2_15min_0[0:0], fa2_15min_0[3:3], fa2_15min_0[5:5]);
  INV I355 (simp2421_0[1:1], fa2_15min_0[6:6]);
  NAND2 I356 (o_0r0[15:15], simp2421_0[0:0], simp2421_0[1:1]);
  NOR3 I357 (simp2431_0[0:0], fa2_15min_0[1:1], fa2_15min_0[2:2], fa2_15min_0[4:4]);
  INV I358 (simp2431_0[1:1], fa2_15min_0[7:7]);
  NAND2 I359 (o_0r1[15:15], simp2431_0[0:0], simp2431_0[1:1]);
  AO222 I360 (ct2__0[15:15], termt_1[15:15], i_0r0[15:15], termt_1[15:15], ct2__0[14:14], i_0r0[15:15], ct2__0[14:14]);
  AO222 I361 (cf2__0[15:15], termf_1[15:15], i_0r1[15:15], termf_1[15:15], cf2__0[14:14], i_0r1[15:15], cf2__0[14:14]);
  C3 I362 (fa2_16min_0[0:0], cf2__0[15:15], i_0r1[16:16], termf_1[16:16]);
  C3 I363 (fa2_16min_0[1:1], cf2__0[15:15], i_0r1[16:16], termt_1[16:16]);
  C3 I364 (fa2_16min_0[2:2], cf2__0[15:15], i_0r0[16:16], termf_1[16:16]);
  C3 I365 (fa2_16min_0[3:3], cf2__0[15:15], i_0r0[16:16], termt_1[16:16]);
  C3 I366 (fa2_16min_0[4:4], ct2__0[15:15], i_0r1[16:16], termf_1[16:16]);
  C3 I367 (fa2_16min_0[5:5], ct2__0[15:15], i_0r1[16:16], termt_1[16:16]);
  C3 I368 (fa2_16min_0[6:6], ct2__0[15:15], i_0r0[16:16], termf_1[16:16]);
  C3 I369 (fa2_16min_0[7:7], ct2__0[15:15], i_0r0[16:16], termt_1[16:16]);
  NOR3 I370 (simp2551_0[0:0], fa2_16min_0[0:0], fa2_16min_0[3:3], fa2_16min_0[5:5]);
  INV I371 (simp2551_0[1:1], fa2_16min_0[6:6]);
  NAND2 I372 (o_0r0[16:16], simp2551_0[0:0], simp2551_0[1:1]);
  NOR3 I373 (simp2561_0[0:0], fa2_16min_0[1:1], fa2_16min_0[2:2], fa2_16min_0[4:4]);
  INV I374 (simp2561_0[1:1], fa2_16min_0[7:7]);
  NAND2 I375 (o_0r1[16:16], simp2561_0[0:0], simp2561_0[1:1]);
  AO222 I376 (ct2__0[16:16], termt_1[16:16], i_0r0[16:16], termt_1[16:16], ct2__0[15:15], i_0r0[16:16], ct2__0[15:15]);
  AO222 I377 (cf2__0[16:16], termf_1[16:16], i_0r1[16:16], termf_1[16:16], cf2__0[15:15], i_0r1[16:16], cf2__0[15:15]);
  C3 I378 (fa2_17min_0[0:0], cf2__0[16:16], i_0r1[17:17], termf_1[17:17]);
  C3 I379 (fa2_17min_0[1:1], cf2__0[16:16], i_0r1[17:17], termt_1[17:17]);
  C3 I380 (fa2_17min_0[2:2], cf2__0[16:16], i_0r0[17:17], termf_1[17:17]);
  C3 I381 (fa2_17min_0[3:3], cf2__0[16:16], i_0r0[17:17], termt_1[17:17]);
  C3 I382 (fa2_17min_0[4:4], ct2__0[16:16], i_0r1[17:17], termf_1[17:17]);
  C3 I383 (fa2_17min_0[5:5], ct2__0[16:16], i_0r1[17:17], termt_1[17:17]);
  C3 I384 (fa2_17min_0[6:6], ct2__0[16:16], i_0r0[17:17], termf_1[17:17]);
  C3 I385 (fa2_17min_0[7:7], ct2__0[16:16], i_0r0[17:17], termt_1[17:17]);
  NOR3 I386 (simp2681_0[0:0], fa2_17min_0[0:0], fa2_17min_0[3:3], fa2_17min_0[5:5]);
  INV I387 (simp2681_0[1:1], fa2_17min_0[6:6]);
  NAND2 I388 (o_0r0[17:17], simp2681_0[0:0], simp2681_0[1:1]);
  NOR3 I389 (simp2691_0[0:0], fa2_17min_0[1:1], fa2_17min_0[2:2], fa2_17min_0[4:4]);
  INV I390 (simp2691_0[1:1], fa2_17min_0[7:7]);
  NAND2 I391 (o_0r1[17:17], simp2691_0[0:0], simp2691_0[1:1]);
  AO222 I392 (ct2__0[17:17], termt_1[17:17], i_0r0[17:17], termt_1[17:17], ct2__0[16:16], i_0r0[17:17], ct2__0[16:16]);
  AO222 I393 (cf2__0[17:17], termf_1[17:17], i_0r1[17:17], termf_1[17:17], cf2__0[16:16], i_0r1[17:17], cf2__0[16:16]);
  C3 I394 (fa2_18min_0[0:0], cf2__0[17:17], i_0r1[18:18], termf_1[18:18]);
  C3 I395 (fa2_18min_0[1:1], cf2__0[17:17], i_0r1[18:18], termt_1[18:18]);
  C3 I396 (fa2_18min_0[2:2], cf2__0[17:17], i_0r0[18:18], termf_1[18:18]);
  C3 I397 (fa2_18min_0[3:3], cf2__0[17:17], i_0r0[18:18], termt_1[18:18]);
  C3 I398 (fa2_18min_0[4:4], ct2__0[17:17], i_0r1[18:18], termf_1[18:18]);
  C3 I399 (fa2_18min_0[5:5], ct2__0[17:17], i_0r1[18:18], termt_1[18:18]);
  C3 I400 (fa2_18min_0[6:6], ct2__0[17:17], i_0r0[18:18], termf_1[18:18]);
  C3 I401 (fa2_18min_0[7:7], ct2__0[17:17], i_0r0[18:18], termt_1[18:18]);
  NOR3 I402 (simp2811_0[0:0], fa2_18min_0[0:0], fa2_18min_0[3:3], fa2_18min_0[5:5]);
  INV I403 (simp2811_0[1:1], fa2_18min_0[6:6]);
  NAND2 I404 (o_0r0[18:18], simp2811_0[0:0], simp2811_0[1:1]);
  NOR3 I405 (simp2821_0[0:0], fa2_18min_0[1:1], fa2_18min_0[2:2], fa2_18min_0[4:4]);
  INV I406 (simp2821_0[1:1], fa2_18min_0[7:7]);
  NAND2 I407 (o_0r1[18:18], simp2821_0[0:0], simp2821_0[1:1]);
  AO222 I408 (ct2__0[18:18], termt_1[18:18], i_0r0[18:18], termt_1[18:18], ct2__0[17:17], i_0r0[18:18], ct2__0[17:17]);
  AO222 I409 (cf2__0[18:18], termf_1[18:18], i_0r1[18:18], termf_1[18:18], cf2__0[17:17], i_0r1[18:18], cf2__0[17:17]);
  C3 I410 (fa2_19min_0[0:0], cf2__0[18:18], i_0r1[19:19], termf_1[19:19]);
  C3 I411 (fa2_19min_0[1:1], cf2__0[18:18], i_0r1[19:19], termt_1[19:19]);
  C3 I412 (fa2_19min_0[2:2], cf2__0[18:18], i_0r0[19:19], termf_1[19:19]);
  C3 I413 (fa2_19min_0[3:3], cf2__0[18:18], i_0r0[19:19], termt_1[19:19]);
  C3 I414 (fa2_19min_0[4:4], ct2__0[18:18], i_0r1[19:19], termf_1[19:19]);
  C3 I415 (fa2_19min_0[5:5], ct2__0[18:18], i_0r1[19:19], termt_1[19:19]);
  C3 I416 (fa2_19min_0[6:6], ct2__0[18:18], i_0r0[19:19], termf_1[19:19]);
  C3 I417 (fa2_19min_0[7:7], ct2__0[18:18], i_0r0[19:19], termt_1[19:19]);
  NOR3 I418 (simp2941_0[0:0], fa2_19min_0[0:0], fa2_19min_0[3:3], fa2_19min_0[5:5]);
  INV I419 (simp2941_0[1:1], fa2_19min_0[6:6]);
  NAND2 I420 (o_0r0[19:19], simp2941_0[0:0], simp2941_0[1:1]);
  NOR3 I421 (simp2951_0[0:0], fa2_19min_0[1:1], fa2_19min_0[2:2], fa2_19min_0[4:4]);
  INV I422 (simp2951_0[1:1], fa2_19min_0[7:7]);
  NAND2 I423 (o_0r1[19:19], simp2951_0[0:0], simp2951_0[1:1]);
  AO222 I424 (ct2__0[19:19], termt_1[19:19], i_0r0[19:19], termt_1[19:19], ct2__0[18:18], i_0r0[19:19], ct2__0[18:18]);
  AO222 I425 (cf2__0[19:19], termf_1[19:19], i_0r1[19:19], termf_1[19:19], cf2__0[18:18], i_0r1[19:19], cf2__0[18:18]);
  C3 I426 (fa2_20min_0[0:0], cf2__0[19:19], i_0r1[20:20], termf_1[20:20]);
  C3 I427 (fa2_20min_0[1:1], cf2__0[19:19], i_0r1[20:20], termt_1[20:20]);
  C3 I428 (fa2_20min_0[2:2], cf2__0[19:19], i_0r0[20:20], termf_1[20:20]);
  C3 I429 (fa2_20min_0[3:3], cf2__0[19:19], i_0r0[20:20], termt_1[20:20]);
  C3 I430 (fa2_20min_0[4:4], ct2__0[19:19], i_0r1[20:20], termf_1[20:20]);
  C3 I431 (fa2_20min_0[5:5], ct2__0[19:19], i_0r1[20:20], termt_1[20:20]);
  C3 I432 (fa2_20min_0[6:6], ct2__0[19:19], i_0r0[20:20], termf_1[20:20]);
  C3 I433 (fa2_20min_0[7:7], ct2__0[19:19], i_0r0[20:20], termt_1[20:20]);
  NOR3 I434 (simp3071_0[0:0], fa2_20min_0[0:0], fa2_20min_0[3:3], fa2_20min_0[5:5]);
  INV I435 (simp3071_0[1:1], fa2_20min_0[6:6]);
  NAND2 I436 (o_0r0[20:20], simp3071_0[0:0], simp3071_0[1:1]);
  NOR3 I437 (simp3081_0[0:0], fa2_20min_0[1:1], fa2_20min_0[2:2], fa2_20min_0[4:4]);
  INV I438 (simp3081_0[1:1], fa2_20min_0[7:7]);
  NAND2 I439 (o_0r1[20:20], simp3081_0[0:0], simp3081_0[1:1]);
  AO222 I440 (ct2__0[20:20], termt_1[20:20], i_0r0[20:20], termt_1[20:20], ct2__0[19:19], i_0r0[20:20], ct2__0[19:19]);
  AO222 I441 (cf2__0[20:20], termf_1[20:20], i_0r1[20:20], termf_1[20:20], cf2__0[19:19], i_0r1[20:20], cf2__0[19:19]);
  C3 I442 (fa2_21min_0[0:0], cf2__0[20:20], i_0r1[21:21], termf_1[21:21]);
  C3 I443 (fa2_21min_0[1:1], cf2__0[20:20], i_0r1[21:21], termt_1[21:21]);
  C3 I444 (fa2_21min_0[2:2], cf2__0[20:20], i_0r0[21:21], termf_1[21:21]);
  C3 I445 (fa2_21min_0[3:3], cf2__0[20:20], i_0r0[21:21], termt_1[21:21]);
  C3 I446 (fa2_21min_0[4:4], ct2__0[20:20], i_0r1[21:21], termf_1[21:21]);
  C3 I447 (fa2_21min_0[5:5], ct2__0[20:20], i_0r1[21:21], termt_1[21:21]);
  C3 I448 (fa2_21min_0[6:6], ct2__0[20:20], i_0r0[21:21], termf_1[21:21]);
  C3 I449 (fa2_21min_0[7:7], ct2__0[20:20], i_0r0[21:21], termt_1[21:21]);
  NOR3 I450 (simp3201_0[0:0], fa2_21min_0[0:0], fa2_21min_0[3:3], fa2_21min_0[5:5]);
  INV I451 (simp3201_0[1:1], fa2_21min_0[6:6]);
  NAND2 I452 (o_0r0[21:21], simp3201_0[0:0], simp3201_0[1:1]);
  NOR3 I453 (simp3211_0[0:0], fa2_21min_0[1:1], fa2_21min_0[2:2], fa2_21min_0[4:4]);
  INV I454 (simp3211_0[1:1], fa2_21min_0[7:7]);
  NAND2 I455 (o_0r1[21:21], simp3211_0[0:0], simp3211_0[1:1]);
  AO222 I456 (ct2__0[21:21], termt_1[21:21], i_0r0[21:21], termt_1[21:21], ct2__0[20:20], i_0r0[21:21], ct2__0[20:20]);
  AO222 I457 (cf2__0[21:21], termf_1[21:21], i_0r1[21:21], termf_1[21:21], cf2__0[20:20], i_0r1[21:21], cf2__0[20:20]);
  C3 I458 (fa2_22min_0[0:0], cf2__0[21:21], i_0r1[22:22], termf_1[22:22]);
  C3 I459 (fa2_22min_0[1:1], cf2__0[21:21], i_0r1[22:22], termt_1[22:22]);
  C3 I460 (fa2_22min_0[2:2], cf2__0[21:21], i_0r0[22:22], termf_1[22:22]);
  C3 I461 (fa2_22min_0[3:3], cf2__0[21:21], i_0r0[22:22], termt_1[22:22]);
  C3 I462 (fa2_22min_0[4:4], ct2__0[21:21], i_0r1[22:22], termf_1[22:22]);
  C3 I463 (fa2_22min_0[5:5], ct2__0[21:21], i_0r1[22:22], termt_1[22:22]);
  C3 I464 (fa2_22min_0[6:6], ct2__0[21:21], i_0r0[22:22], termf_1[22:22]);
  C3 I465 (fa2_22min_0[7:7], ct2__0[21:21], i_0r0[22:22], termt_1[22:22]);
  NOR3 I466 (simp3331_0[0:0], fa2_22min_0[0:0], fa2_22min_0[3:3], fa2_22min_0[5:5]);
  INV I467 (simp3331_0[1:1], fa2_22min_0[6:6]);
  NAND2 I468 (o_0r0[22:22], simp3331_0[0:0], simp3331_0[1:1]);
  NOR3 I469 (simp3341_0[0:0], fa2_22min_0[1:1], fa2_22min_0[2:2], fa2_22min_0[4:4]);
  INV I470 (simp3341_0[1:1], fa2_22min_0[7:7]);
  NAND2 I471 (o_0r1[22:22], simp3341_0[0:0], simp3341_0[1:1]);
  AO222 I472 (ct2__0[22:22], termt_1[22:22], i_0r0[22:22], termt_1[22:22], ct2__0[21:21], i_0r0[22:22], ct2__0[21:21]);
  AO222 I473 (cf2__0[22:22], termf_1[22:22], i_0r1[22:22], termf_1[22:22], cf2__0[21:21], i_0r1[22:22], cf2__0[21:21]);
  C3 I474 (fa2_23min_0[0:0], cf2__0[22:22], i_0r1[23:23], termf_1[23:23]);
  C3 I475 (fa2_23min_0[1:1], cf2__0[22:22], i_0r1[23:23], termt_1[23:23]);
  C3 I476 (fa2_23min_0[2:2], cf2__0[22:22], i_0r0[23:23], termf_1[23:23]);
  C3 I477 (fa2_23min_0[3:3], cf2__0[22:22], i_0r0[23:23], termt_1[23:23]);
  C3 I478 (fa2_23min_0[4:4], ct2__0[22:22], i_0r1[23:23], termf_1[23:23]);
  C3 I479 (fa2_23min_0[5:5], ct2__0[22:22], i_0r1[23:23], termt_1[23:23]);
  C3 I480 (fa2_23min_0[6:6], ct2__0[22:22], i_0r0[23:23], termf_1[23:23]);
  C3 I481 (fa2_23min_0[7:7], ct2__0[22:22], i_0r0[23:23], termt_1[23:23]);
  NOR3 I482 (simp3461_0[0:0], fa2_23min_0[0:0], fa2_23min_0[3:3], fa2_23min_0[5:5]);
  INV I483 (simp3461_0[1:1], fa2_23min_0[6:6]);
  NAND2 I484 (o_0r0[23:23], simp3461_0[0:0], simp3461_0[1:1]);
  NOR3 I485 (simp3471_0[0:0], fa2_23min_0[1:1], fa2_23min_0[2:2], fa2_23min_0[4:4]);
  INV I486 (simp3471_0[1:1], fa2_23min_0[7:7]);
  NAND2 I487 (o_0r1[23:23], simp3471_0[0:0], simp3471_0[1:1]);
  AO222 I488 (ct2__0[23:23], termt_1[23:23], i_0r0[23:23], termt_1[23:23], ct2__0[22:22], i_0r0[23:23], ct2__0[22:22]);
  AO222 I489 (cf2__0[23:23], termf_1[23:23], i_0r1[23:23], termf_1[23:23], cf2__0[22:22], i_0r1[23:23], cf2__0[22:22]);
  C3 I490 (fa2_24min_0[0:0], cf2__0[23:23], i_0r1[24:24], termf_1[24:24]);
  C3 I491 (fa2_24min_0[1:1], cf2__0[23:23], i_0r1[24:24], termt_1[24:24]);
  C3 I492 (fa2_24min_0[2:2], cf2__0[23:23], i_0r0[24:24], termf_1[24:24]);
  C3 I493 (fa2_24min_0[3:3], cf2__0[23:23], i_0r0[24:24], termt_1[24:24]);
  C3 I494 (fa2_24min_0[4:4], ct2__0[23:23], i_0r1[24:24], termf_1[24:24]);
  C3 I495 (fa2_24min_0[5:5], ct2__0[23:23], i_0r1[24:24], termt_1[24:24]);
  C3 I496 (fa2_24min_0[6:6], ct2__0[23:23], i_0r0[24:24], termf_1[24:24]);
  C3 I497 (fa2_24min_0[7:7], ct2__0[23:23], i_0r0[24:24], termt_1[24:24]);
  NOR3 I498 (simp3591_0[0:0], fa2_24min_0[0:0], fa2_24min_0[3:3], fa2_24min_0[5:5]);
  INV I499 (simp3591_0[1:1], fa2_24min_0[6:6]);
  NAND2 I500 (o_0r0[24:24], simp3591_0[0:0], simp3591_0[1:1]);
  NOR3 I501 (simp3601_0[0:0], fa2_24min_0[1:1], fa2_24min_0[2:2], fa2_24min_0[4:4]);
  INV I502 (simp3601_0[1:1], fa2_24min_0[7:7]);
  NAND2 I503 (o_0r1[24:24], simp3601_0[0:0], simp3601_0[1:1]);
  AO222 I504 (ct2__0[24:24], termt_1[24:24], i_0r0[24:24], termt_1[24:24], ct2__0[23:23], i_0r0[24:24], ct2__0[23:23]);
  AO222 I505 (cf2__0[24:24], termf_1[24:24], i_0r1[24:24], termf_1[24:24], cf2__0[23:23], i_0r1[24:24], cf2__0[23:23]);
  C3 I506 (fa2_25min_0[0:0], cf2__0[24:24], i_0r1[25:25], termf_1[25:25]);
  C3 I507 (fa2_25min_0[1:1], cf2__0[24:24], i_0r1[25:25], termt_1[25:25]);
  C3 I508 (fa2_25min_0[2:2], cf2__0[24:24], i_0r0[25:25], termf_1[25:25]);
  C3 I509 (fa2_25min_0[3:3], cf2__0[24:24], i_0r0[25:25], termt_1[25:25]);
  C3 I510 (fa2_25min_0[4:4], ct2__0[24:24], i_0r1[25:25], termf_1[25:25]);
  C3 I511 (fa2_25min_0[5:5], ct2__0[24:24], i_0r1[25:25], termt_1[25:25]);
  C3 I512 (fa2_25min_0[6:6], ct2__0[24:24], i_0r0[25:25], termf_1[25:25]);
  C3 I513 (fa2_25min_0[7:7], ct2__0[24:24], i_0r0[25:25], termt_1[25:25]);
  NOR3 I514 (simp3721_0[0:0], fa2_25min_0[0:0], fa2_25min_0[3:3], fa2_25min_0[5:5]);
  INV I515 (simp3721_0[1:1], fa2_25min_0[6:6]);
  NAND2 I516 (o_0r0[25:25], simp3721_0[0:0], simp3721_0[1:1]);
  NOR3 I517 (simp3731_0[0:0], fa2_25min_0[1:1], fa2_25min_0[2:2], fa2_25min_0[4:4]);
  INV I518 (simp3731_0[1:1], fa2_25min_0[7:7]);
  NAND2 I519 (o_0r1[25:25], simp3731_0[0:0], simp3731_0[1:1]);
  AO222 I520 (ct2__0[25:25], termt_1[25:25], i_0r0[25:25], termt_1[25:25], ct2__0[24:24], i_0r0[25:25], ct2__0[24:24]);
  AO222 I521 (cf2__0[25:25], termf_1[25:25], i_0r1[25:25], termf_1[25:25], cf2__0[24:24], i_0r1[25:25], cf2__0[24:24]);
  C3 I522 (fa2_26min_0[0:0], cf2__0[25:25], i_0r1[26:26], termf_1[26:26]);
  C3 I523 (fa2_26min_0[1:1], cf2__0[25:25], i_0r1[26:26], termt_1[26:26]);
  C3 I524 (fa2_26min_0[2:2], cf2__0[25:25], i_0r0[26:26], termf_1[26:26]);
  C3 I525 (fa2_26min_0[3:3], cf2__0[25:25], i_0r0[26:26], termt_1[26:26]);
  C3 I526 (fa2_26min_0[4:4], ct2__0[25:25], i_0r1[26:26], termf_1[26:26]);
  C3 I527 (fa2_26min_0[5:5], ct2__0[25:25], i_0r1[26:26], termt_1[26:26]);
  C3 I528 (fa2_26min_0[6:6], ct2__0[25:25], i_0r0[26:26], termf_1[26:26]);
  C3 I529 (fa2_26min_0[7:7], ct2__0[25:25], i_0r0[26:26], termt_1[26:26]);
  NOR3 I530 (simp3851_0[0:0], fa2_26min_0[0:0], fa2_26min_0[3:3], fa2_26min_0[5:5]);
  INV I531 (simp3851_0[1:1], fa2_26min_0[6:6]);
  NAND2 I532 (o_0r0[26:26], simp3851_0[0:0], simp3851_0[1:1]);
  NOR3 I533 (simp3861_0[0:0], fa2_26min_0[1:1], fa2_26min_0[2:2], fa2_26min_0[4:4]);
  INV I534 (simp3861_0[1:1], fa2_26min_0[7:7]);
  NAND2 I535 (o_0r1[26:26], simp3861_0[0:0], simp3861_0[1:1]);
  AO222 I536 (ct2__0[26:26], termt_1[26:26], i_0r0[26:26], termt_1[26:26], ct2__0[25:25], i_0r0[26:26], ct2__0[25:25]);
  AO222 I537 (cf2__0[26:26], termf_1[26:26], i_0r1[26:26], termf_1[26:26], cf2__0[25:25], i_0r1[26:26], cf2__0[25:25]);
  C3 I538 (fa2_27min_0[0:0], cf2__0[26:26], i_0r1[27:27], termf_1[27:27]);
  C3 I539 (fa2_27min_0[1:1], cf2__0[26:26], i_0r1[27:27], termt_1[27:27]);
  C3 I540 (fa2_27min_0[2:2], cf2__0[26:26], i_0r0[27:27], termf_1[27:27]);
  C3 I541 (fa2_27min_0[3:3], cf2__0[26:26], i_0r0[27:27], termt_1[27:27]);
  C3 I542 (fa2_27min_0[4:4], ct2__0[26:26], i_0r1[27:27], termf_1[27:27]);
  C3 I543 (fa2_27min_0[5:5], ct2__0[26:26], i_0r1[27:27], termt_1[27:27]);
  C3 I544 (fa2_27min_0[6:6], ct2__0[26:26], i_0r0[27:27], termf_1[27:27]);
  C3 I545 (fa2_27min_0[7:7], ct2__0[26:26], i_0r0[27:27], termt_1[27:27]);
  NOR3 I546 (simp3981_0[0:0], fa2_27min_0[0:0], fa2_27min_0[3:3], fa2_27min_0[5:5]);
  INV I547 (simp3981_0[1:1], fa2_27min_0[6:6]);
  NAND2 I548 (o_0r0[27:27], simp3981_0[0:0], simp3981_0[1:1]);
  NOR3 I549 (simp3991_0[0:0], fa2_27min_0[1:1], fa2_27min_0[2:2], fa2_27min_0[4:4]);
  INV I550 (simp3991_0[1:1], fa2_27min_0[7:7]);
  NAND2 I551 (o_0r1[27:27], simp3991_0[0:0], simp3991_0[1:1]);
  AO222 I552 (ct2__0[27:27], termt_1[27:27], i_0r0[27:27], termt_1[27:27], ct2__0[26:26], i_0r0[27:27], ct2__0[26:26]);
  AO222 I553 (cf2__0[27:27], termf_1[27:27], i_0r1[27:27], termf_1[27:27], cf2__0[26:26], i_0r1[27:27], cf2__0[26:26]);
  C3 I554 (fa2_28min_0[0:0], cf2__0[27:27], i_0r1[28:28], termf_1[28:28]);
  C3 I555 (fa2_28min_0[1:1], cf2__0[27:27], i_0r1[28:28], termt_1[28:28]);
  C3 I556 (fa2_28min_0[2:2], cf2__0[27:27], i_0r0[28:28], termf_1[28:28]);
  C3 I557 (fa2_28min_0[3:3], cf2__0[27:27], i_0r0[28:28], termt_1[28:28]);
  C3 I558 (fa2_28min_0[4:4], ct2__0[27:27], i_0r1[28:28], termf_1[28:28]);
  C3 I559 (fa2_28min_0[5:5], ct2__0[27:27], i_0r1[28:28], termt_1[28:28]);
  C3 I560 (fa2_28min_0[6:6], ct2__0[27:27], i_0r0[28:28], termf_1[28:28]);
  C3 I561 (fa2_28min_0[7:7], ct2__0[27:27], i_0r0[28:28], termt_1[28:28]);
  NOR3 I562 (simp4111_0[0:0], fa2_28min_0[0:0], fa2_28min_0[3:3], fa2_28min_0[5:5]);
  INV I563 (simp4111_0[1:1], fa2_28min_0[6:6]);
  NAND2 I564 (o_0r0[28:28], simp4111_0[0:0], simp4111_0[1:1]);
  NOR3 I565 (simp4121_0[0:0], fa2_28min_0[1:1], fa2_28min_0[2:2], fa2_28min_0[4:4]);
  INV I566 (simp4121_0[1:1], fa2_28min_0[7:7]);
  NAND2 I567 (o_0r1[28:28], simp4121_0[0:0], simp4121_0[1:1]);
  AO222 I568 (ct2__0[28:28], termt_1[28:28], i_0r0[28:28], termt_1[28:28], ct2__0[27:27], i_0r0[28:28], ct2__0[27:27]);
  AO222 I569 (cf2__0[28:28], termf_1[28:28], i_0r1[28:28], termf_1[28:28], cf2__0[27:27], i_0r1[28:28], cf2__0[27:27]);
  C3 I570 (fa2_29min_0[0:0], cf2__0[28:28], i_0r1[29:29], termf_1[29:29]);
  C3 I571 (fa2_29min_0[1:1], cf2__0[28:28], i_0r1[29:29], termt_1[29:29]);
  C3 I572 (fa2_29min_0[2:2], cf2__0[28:28], i_0r0[29:29], termf_1[29:29]);
  C3 I573 (fa2_29min_0[3:3], cf2__0[28:28], i_0r0[29:29], termt_1[29:29]);
  C3 I574 (fa2_29min_0[4:4], ct2__0[28:28], i_0r1[29:29], termf_1[29:29]);
  C3 I575 (fa2_29min_0[5:5], ct2__0[28:28], i_0r1[29:29], termt_1[29:29]);
  C3 I576 (fa2_29min_0[6:6], ct2__0[28:28], i_0r0[29:29], termf_1[29:29]);
  C3 I577 (fa2_29min_0[7:7], ct2__0[28:28], i_0r0[29:29], termt_1[29:29]);
  NOR3 I578 (simp4241_0[0:0], fa2_29min_0[0:0], fa2_29min_0[3:3], fa2_29min_0[5:5]);
  INV I579 (simp4241_0[1:1], fa2_29min_0[6:6]);
  NAND2 I580 (o_0r0[29:29], simp4241_0[0:0], simp4241_0[1:1]);
  NOR3 I581 (simp4251_0[0:0], fa2_29min_0[1:1], fa2_29min_0[2:2], fa2_29min_0[4:4]);
  INV I582 (simp4251_0[1:1], fa2_29min_0[7:7]);
  NAND2 I583 (o_0r1[29:29], simp4251_0[0:0], simp4251_0[1:1]);
  AO222 I584 (ct2__0[29:29], termt_1[29:29], i_0r0[29:29], termt_1[29:29], ct2__0[28:28], i_0r0[29:29], ct2__0[28:28]);
  AO222 I585 (cf2__0[29:29], termf_1[29:29], i_0r1[29:29], termf_1[29:29], cf2__0[28:28], i_0r1[29:29], cf2__0[28:28]);
  C3 I586 (fa2_30min_0[0:0], cf2__0[29:29], i_0r1[30:30], termf_1[30:30]);
  C3 I587 (fa2_30min_0[1:1], cf2__0[29:29], i_0r1[30:30], termt_1[30:30]);
  C3 I588 (fa2_30min_0[2:2], cf2__0[29:29], i_0r0[30:30], termf_1[30:30]);
  C3 I589 (fa2_30min_0[3:3], cf2__0[29:29], i_0r0[30:30], termt_1[30:30]);
  C3 I590 (fa2_30min_0[4:4], ct2__0[29:29], i_0r1[30:30], termf_1[30:30]);
  C3 I591 (fa2_30min_0[5:5], ct2__0[29:29], i_0r1[30:30], termt_1[30:30]);
  C3 I592 (fa2_30min_0[6:6], ct2__0[29:29], i_0r0[30:30], termf_1[30:30]);
  C3 I593 (fa2_30min_0[7:7], ct2__0[29:29], i_0r0[30:30], termt_1[30:30]);
  NOR3 I594 (simp4371_0[0:0], fa2_30min_0[0:0], fa2_30min_0[3:3], fa2_30min_0[5:5]);
  INV I595 (simp4371_0[1:1], fa2_30min_0[6:6]);
  NAND2 I596 (o_0r0[30:30], simp4371_0[0:0], simp4371_0[1:1]);
  NOR3 I597 (simp4381_0[0:0], fa2_30min_0[1:1], fa2_30min_0[2:2], fa2_30min_0[4:4]);
  INV I598 (simp4381_0[1:1], fa2_30min_0[7:7]);
  NAND2 I599 (o_0r1[30:30], simp4381_0[0:0], simp4381_0[1:1]);
  AO222 I600 (ct2__0[30:30], termt_1[30:30], i_0r0[30:30], termt_1[30:30], ct2__0[29:29], i_0r0[30:30], ct2__0[29:29]);
  AO222 I601 (cf2__0[30:30], termf_1[30:30], i_0r1[30:30], termf_1[30:30], cf2__0[29:29], i_0r1[30:30], cf2__0[29:29]);
  C3 I602 (fa2_31min_0[0:0], cf2__0[30:30], i_0r1[31:31], termf_1[31:31]);
  C3 I603 (fa2_31min_0[1:1], cf2__0[30:30], i_0r1[31:31], termt_1[31:31]);
  C3 I604 (fa2_31min_0[2:2], cf2__0[30:30], i_0r0[31:31], termf_1[31:31]);
  C3 I605 (fa2_31min_0[3:3], cf2__0[30:30], i_0r0[31:31], termt_1[31:31]);
  C3 I606 (fa2_31min_0[4:4], ct2__0[30:30], i_0r1[31:31], termf_1[31:31]);
  C3 I607 (fa2_31min_0[5:5], ct2__0[30:30], i_0r1[31:31], termt_1[31:31]);
  C3 I608 (fa2_31min_0[6:6], ct2__0[30:30], i_0r0[31:31], termf_1[31:31]);
  C3 I609 (fa2_31min_0[7:7], ct2__0[30:30], i_0r0[31:31], termt_1[31:31]);
  NOR3 I610 (simp4501_0[0:0], fa2_31min_0[0:0], fa2_31min_0[3:3], fa2_31min_0[5:5]);
  INV I611 (simp4501_0[1:1], fa2_31min_0[6:6]);
  NAND2 I612 (o_0r0[31:31], simp4501_0[0:0], simp4501_0[1:1]);
  NOR3 I613 (simp4511_0[0:0], fa2_31min_0[1:1], fa2_31min_0[2:2], fa2_31min_0[4:4]);
  INV I614 (simp4511_0[1:1], fa2_31min_0[7:7]);
  NAND2 I615 (o_0r1[31:31], simp4511_0[0:0], simp4511_0[1:1]);
  AO222 I616 (ct2__0[31:31], termt_1[31:31], i_0r0[31:31], termt_1[31:31], ct2__0[30:30], i_0r0[31:31], ct2__0[30:30]);
  AO222 I617 (cf2__0[31:31], termf_1[31:31], i_0r1[31:31], termf_1[31:31], cf2__0[30:30], i_0r1[31:31], cf2__0[30:30]);
  BUFF I618 (i_0a, o_0a);
endmodule

// tkf4mo0w0_o0w3 TeakF [0,0] [One 4,Many [0,3]]
module tkf4mo0w0_o0w3 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [2:0] o_1r0;
  output [2:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire comp_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0, i_0r0[3:3], i_0r1[3:3]);
  BUFF I2 (ucomplete_0, comp_0);
  C2 I3 (acomplete_0, ucomplete_0, icomplete_0);
  C2 I4 (o_1r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I5 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I6 (o_1r0[2:2], i_0r0[2:2]);
  C2 I7 (o_1r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I8 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I9 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I10 (o_0r, icomplete_0);
  C3 I11 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tks1_o0w1_0o0w0_1o0w0 TeakS (0+:1) [([Imp 0 0],0),([Imp 1 0],0)] [One 1,Many [0,0]]
module tks1_o0w1_0o0w0_1o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire comp_0;
  BUFF I0 (sel_0, match0_0);
  BUFF I1 (match0_0, i_0r0);
  BUFF I2 (sel_1, match1_0);
  BUFF I3 (match1_0, i_0r1);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0, i_0r0, i_0r1);
  BUFF I7 (icomplete_0, comp_0);
  BUFF I8 (o_0r, gsel_0);
  BUFF I9 (o_1r, gsel_1);
  OR2 I10 (oack_0, o_0a, o_1a);
  C2 I11 (i_0a, oack_0, icomplete_0);
endmodule

// tkm2x0b TeakM [Many [0,0],One 0]
module tkm2x0b (i_0r, i_0a, i_1r, i_1a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  NOR2 I2 (nchosen_0, o_0r, o_0a);
  OR2 I3 (o_0r, choice_0, choice_1);
  C2R I4 (i_0a, choice_0, o_0a, reset);
  C2R I5 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj64m32_32 TeakJ [Many [32,32],One 64]
module tkj64m32_32 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [63:0] o_0r0;
  output [63:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [63:0] joinf_0;
  wire [63:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joinf_0[34:34], i_1r0[2:2]);
  BUFF I35 (joinf_0[35:35], i_1r0[3:3]);
  BUFF I36 (joinf_0[36:36], i_1r0[4:4]);
  BUFF I37 (joinf_0[37:37], i_1r0[5:5]);
  BUFF I38 (joinf_0[38:38], i_1r0[6:6]);
  BUFF I39 (joinf_0[39:39], i_1r0[7:7]);
  BUFF I40 (joinf_0[40:40], i_1r0[8:8]);
  BUFF I41 (joinf_0[41:41], i_1r0[9:9]);
  BUFF I42 (joinf_0[42:42], i_1r0[10:10]);
  BUFF I43 (joinf_0[43:43], i_1r0[11:11]);
  BUFF I44 (joinf_0[44:44], i_1r0[12:12]);
  BUFF I45 (joinf_0[45:45], i_1r0[13:13]);
  BUFF I46 (joinf_0[46:46], i_1r0[14:14]);
  BUFF I47 (joinf_0[47:47], i_1r0[15:15]);
  BUFF I48 (joinf_0[48:48], i_1r0[16:16]);
  BUFF I49 (joinf_0[49:49], i_1r0[17:17]);
  BUFF I50 (joinf_0[50:50], i_1r0[18:18]);
  BUFF I51 (joinf_0[51:51], i_1r0[19:19]);
  BUFF I52 (joinf_0[52:52], i_1r0[20:20]);
  BUFF I53 (joinf_0[53:53], i_1r0[21:21]);
  BUFF I54 (joinf_0[54:54], i_1r0[22:22]);
  BUFF I55 (joinf_0[55:55], i_1r0[23:23]);
  BUFF I56 (joinf_0[56:56], i_1r0[24:24]);
  BUFF I57 (joinf_0[57:57], i_1r0[25:25]);
  BUFF I58 (joinf_0[58:58], i_1r0[26:26]);
  BUFF I59 (joinf_0[59:59], i_1r0[27:27]);
  BUFF I60 (joinf_0[60:60], i_1r0[28:28]);
  BUFF I61 (joinf_0[61:61], i_1r0[29:29]);
  BUFF I62 (joinf_0[62:62], i_1r0[30:30]);
  BUFF I63 (joinf_0[63:63], i_1r0[31:31]);
  BUFF I64 (joint_0[0:0], i_0r1[0:0]);
  BUFF I65 (joint_0[1:1], i_0r1[1:1]);
  BUFF I66 (joint_0[2:2], i_0r1[2:2]);
  BUFF I67 (joint_0[3:3], i_0r1[3:3]);
  BUFF I68 (joint_0[4:4], i_0r1[4:4]);
  BUFF I69 (joint_0[5:5], i_0r1[5:5]);
  BUFF I70 (joint_0[6:6], i_0r1[6:6]);
  BUFF I71 (joint_0[7:7], i_0r1[7:7]);
  BUFF I72 (joint_0[8:8], i_0r1[8:8]);
  BUFF I73 (joint_0[9:9], i_0r1[9:9]);
  BUFF I74 (joint_0[10:10], i_0r1[10:10]);
  BUFF I75 (joint_0[11:11], i_0r1[11:11]);
  BUFF I76 (joint_0[12:12], i_0r1[12:12]);
  BUFF I77 (joint_0[13:13], i_0r1[13:13]);
  BUFF I78 (joint_0[14:14], i_0r1[14:14]);
  BUFF I79 (joint_0[15:15], i_0r1[15:15]);
  BUFF I80 (joint_0[16:16], i_0r1[16:16]);
  BUFF I81 (joint_0[17:17], i_0r1[17:17]);
  BUFF I82 (joint_0[18:18], i_0r1[18:18]);
  BUFF I83 (joint_0[19:19], i_0r1[19:19]);
  BUFF I84 (joint_0[20:20], i_0r1[20:20]);
  BUFF I85 (joint_0[21:21], i_0r1[21:21]);
  BUFF I86 (joint_0[22:22], i_0r1[22:22]);
  BUFF I87 (joint_0[23:23], i_0r1[23:23]);
  BUFF I88 (joint_0[24:24], i_0r1[24:24]);
  BUFF I89 (joint_0[25:25], i_0r1[25:25]);
  BUFF I90 (joint_0[26:26], i_0r1[26:26]);
  BUFF I91 (joint_0[27:27], i_0r1[27:27]);
  BUFF I92 (joint_0[28:28], i_0r1[28:28]);
  BUFF I93 (joint_0[29:29], i_0r1[29:29]);
  BUFF I94 (joint_0[30:30], i_0r1[30:30]);
  BUFF I95 (joint_0[31:31], i_0r1[31:31]);
  BUFF I96 (joint_0[32:32], i_1r1[0:0]);
  BUFF I97 (joint_0[33:33], i_1r1[1:1]);
  BUFF I98 (joint_0[34:34], i_1r1[2:2]);
  BUFF I99 (joint_0[35:35], i_1r1[3:3]);
  BUFF I100 (joint_0[36:36], i_1r1[4:4]);
  BUFF I101 (joint_0[37:37], i_1r1[5:5]);
  BUFF I102 (joint_0[38:38], i_1r1[6:6]);
  BUFF I103 (joint_0[39:39], i_1r1[7:7]);
  BUFF I104 (joint_0[40:40], i_1r1[8:8]);
  BUFF I105 (joint_0[41:41], i_1r1[9:9]);
  BUFF I106 (joint_0[42:42], i_1r1[10:10]);
  BUFF I107 (joint_0[43:43], i_1r1[11:11]);
  BUFF I108 (joint_0[44:44], i_1r1[12:12]);
  BUFF I109 (joint_0[45:45], i_1r1[13:13]);
  BUFF I110 (joint_0[46:46], i_1r1[14:14]);
  BUFF I111 (joint_0[47:47], i_1r1[15:15]);
  BUFF I112 (joint_0[48:48], i_1r1[16:16]);
  BUFF I113 (joint_0[49:49], i_1r1[17:17]);
  BUFF I114 (joint_0[50:50], i_1r1[18:18]);
  BUFF I115 (joint_0[51:51], i_1r1[19:19]);
  BUFF I116 (joint_0[52:52], i_1r1[20:20]);
  BUFF I117 (joint_0[53:53], i_1r1[21:21]);
  BUFF I118 (joint_0[54:54], i_1r1[22:22]);
  BUFF I119 (joint_0[55:55], i_1r1[23:23]);
  BUFF I120 (joint_0[56:56], i_1r1[24:24]);
  BUFF I121 (joint_0[57:57], i_1r1[25:25]);
  BUFF I122 (joint_0[58:58], i_1r1[26:26]);
  BUFF I123 (joint_0[59:59], i_1r1[27:27]);
  BUFF I124 (joint_0[60:60], i_1r1[28:28]);
  BUFF I125 (joint_0[61:61], i_1r1[29:29]);
  BUFF I126 (joint_0[62:62], i_1r1[30:30]);
  BUFF I127 (joint_0[63:63], i_1r1[31:31]);
  OR2 I128 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I129 (icomplete_0, dcomplete_0);
  C2 I130 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I131 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I132 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I133 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I134 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I135 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I136 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I137 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I138 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I139 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I140 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I141 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I142 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I143 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I144 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I145 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I146 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I147 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I148 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I149 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I150 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I151 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I152 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I153 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I154 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I155 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I156 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I157 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I158 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I159 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I160 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I161 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I162 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I163 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I164 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I165 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I166 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I167 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I168 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I169 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I170 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I171 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I172 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I173 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I174 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I175 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I176 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I177 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I178 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I179 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I180 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I181 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I182 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I183 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I184 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I185 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I186 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I187 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I188 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I189 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I190 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I191 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I192 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I193 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I194 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I195 (o_0r1[1:1], joint_0[1:1]);
  BUFF I196 (o_0r1[2:2], joint_0[2:2]);
  BUFF I197 (o_0r1[3:3], joint_0[3:3]);
  BUFF I198 (o_0r1[4:4], joint_0[4:4]);
  BUFF I199 (o_0r1[5:5], joint_0[5:5]);
  BUFF I200 (o_0r1[6:6], joint_0[6:6]);
  BUFF I201 (o_0r1[7:7], joint_0[7:7]);
  BUFF I202 (o_0r1[8:8], joint_0[8:8]);
  BUFF I203 (o_0r1[9:9], joint_0[9:9]);
  BUFF I204 (o_0r1[10:10], joint_0[10:10]);
  BUFF I205 (o_0r1[11:11], joint_0[11:11]);
  BUFF I206 (o_0r1[12:12], joint_0[12:12]);
  BUFF I207 (o_0r1[13:13], joint_0[13:13]);
  BUFF I208 (o_0r1[14:14], joint_0[14:14]);
  BUFF I209 (o_0r1[15:15], joint_0[15:15]);
  BUFF I210 (o_0r1[16:16], joint_0[16:16]);
  BUFF I211 (o_0r1[17:17], joint_0[17:17]);
  BUFF I212 (o_0r1[18:18], joint_0[18:18]);
  BUFF I213 (o_0r1[19:19], joint_0[19:19]);
  BUFF I214 (o_0r1[20:20], joint_0[20:20]);
  BUFF I215 (o_0r1[21:21], joint_0[21:21]);
  BUFF I216 (o_0r1[22:22], joint_0[22:22]);
  BUFF I217 (o_0r1[23:23], joint_0[23:23]);
  BUFF I218 (o_0r1[24:24], joint_0[24:24]);
  BUFF I219 (o_0r1[25:25], joint_0[25:25]);
  BUFF I220 (o_0r1[26:26], joint_0[26:26]);
  BUFF I221 (o_0r1[27:27], joint_0[27:27]);
  BUFF I222 (o_0r1[28:28], joint_0[28:28]);
  BUFF I223 (o_0r1[29:29], joint_0[29:29]);
  BUFF I224 (o_0r1[30:30], joint_0[30:30]);
  BUFF I225 (o_0r1[31:31], joint_0[31:31]);
  BUFF I226 (o_0r1[32:32], joint_0[32:32]);
  BUFF I227 (o_0r1[33:33], joint_0[33:33]);
  BUFF I228 (o_0r1[34:34], joint_0[34:34]);
  BUFF I229 (o_0r1[35:35], joint_0[35:35]);
  BUFF I230 (o_0r1[36:36], joint_0[36:36]);
  BUFF I231 (o_0r1[37:37], joint_0[37:37]);
  BUFF I232 (o_0r1[38:38], joint_0[38:38]);
  BUFF I233 (o_0r1[39:39], joint_0[39:39]);
  BUFF I234 (o_0r1[40:40], joint_0[40:40]);
  BUFF I235 (o_0r1[41:41], joint_0[41:41]);
  BUFF I236 (o_0r1[42:42], joint_0[42:42]);
  BUFF I237 (o_0r1[43:43], joint_0[43:43]);
  BUFF I238 (o_0r1[44:44], joint_0[44:44]);
  BUFF I239 (o_0r1[45:45], joint_0[45:45]);
  BUFF I240 (o_0r1[46:46], joint_0[46:46]);
  BUFF I241 (o_0r1[47:47], joint_0[47:47]);
  BUFF I242 (o_0r1[48:48], joint_0[48:48]);
  BUFF I243 (o_0r1[49:49], joint_0[49:49]);
  BUFF I244 (o_0r1[50:50], joint_0[50:50]);
  BUFF I245 (o_0r1[51:51], joint_0[51:51]);
  BUFF I246 (o_0r1[52:52], joint_0[52:52]);
  BUFF I247 (o_0r1[53:53], joint_0[53:53]);
  BUFF I248 (o_0r1[54:54], joint_0[54:54]);
  BUFF I249 (o_0r1[55:55], joint_0[55:55]);
  BUFF I250 (o_0r1[56:56], joint_0[56:56]);
  BUFF I251 (o_0r1[57:57], joint_0[57:57]);
  BUFF I252 (o_0r1[58:58], joint_0[58:58]);
  BUFF I253 (o_0r1[59:59], joint_0[59:59]);
  BUFF I254 (o_0r1[60:60], joint_0[60:60]);
  BUFF I255 (o_0r1[61:61], joint_0[61:61]);
  BUFF I256 (o_0r1[62:62], joint_0[62:62]);
  BUFF I257 (o_0r1[63:63], joint_0[63:63]);
  BUFF I258 (i_0a, o_0a);
  BUFF I259 (i_1a, o_0a);
endmodule

// tko64m33_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32),(0,31+:1)]),
//     (2,TeakOAppend 1 [(0,32+:32),(0,63+:1)]),
//     (3,TeakOp TeakOpAdd [(1,0+:33),(2,0+:33)])] [One 64,One 33]
module tko64m33_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire [32:0] termf_1;
  wire [32:0] termf_2;
  wire [32:0] termt_1;
  wire [32:0] termt_2;
  wire [32:0] cf3__0;
  wire [32:0] ct3__0;
  wire [3:0] ha3__0;
  wire [7:0] fa3_1min_0;
  wire [1:0] simp1561_0;
  wire [1:0] simp1571_0;
  wire [7:0] fa3_2min_0;
  wire [1:0] simp1691_0;
  wire [1:0] simp1701_0;
  wire [7:0] fa3_3min_0;
  wire [1:0] simp1821_0;
  wire [1:0] simp1831_0;
  wire [7:0] fa3_4min_0;
  wire [1:0] simp1951_0;
  wire [1:0] simp1961_0;
  wire [7:0] fa3_5min_0;
  wire [1:0] simp2081_0;
  wire [1:0] simp2091_0;
  wire [7:0] fa3_6min_0;
  wire [1:0] simp2211_0;
  wire [1:0] simp2221_0;
  wire [7:0] fa3_7min_0;
  wire [1:0] simp2341_0;
  wire [1:0] simp2351_0;
  wire [7:0] fa3_8min_0;
  wire [1:0] simp2471_0;
  wire [1:0] simp2481_0;
  wire [7:0] fa3_9min_0;
  wire [1:0] simp2601_0;
  wire [1:0] simp2611_0;
  wire [7:0] fa3_10min_0;
  wire [1:0] simp2731_0;
  wire [1:0] simp2741_0;
  wire [7:0] fa3_11min_0;
  wire [1:0] simp2861_0;
  wire [1:0] simp2871_0;
  wire [7:0] fa3_12min_0;
  wire [1:0] simp2991_0;
  wire [1:0] simp3001_0;
  wire [7:0] fa3_13min_0;
  wire [1:0] simp3121_0;
  wire [1:0] simp3131_0;
  wire [7:0] fa3_14min_0;
  wire [1:0] simp3251_0;
  wire [1:0] simp3261_0;
  wire [7:0] fa3_15min_0;
  wire [1:0] simp3381_0;
  wire [1:0] simp3391_0;
  wire [7:0] fa3_16min_0;
  wire [1:0] simp3511_0;
  wire [1:0] simp3521_0;
  wire [7:0] fa3_17min_0;
  wire [1:0] simp3641_0;
  wire [1:0] simp3651_0;
  wire [7:0] fa3_18min_0;
  wire [1:0] simp3771_0;
  wire [1:0] simp3781_0;
  wire [7:0] fa3_19min_0;
  wire [1:0] simp3901_0;
  wire [1:0] simp3911_0;
  wire [7:0] fa3_20min_0;
  wire [1:0] simp4031_0;
  wire [1:0] simp4041_0;
  wire [7:0] fa3_21min_0;
  wire [1:0] simp4161_0;
  wire [1:0] simp4171_0;
  wire [7:0] fa3_22min_0;
  wire [1:0] simp4291_0;
  wire [1:0] simp4301_0;
  wire [7:0] fa3_23min_0;
  wire [1:0] simp4421_0;
  wire [1:0] simp4431_0;
  wire [7:0] fa3_24min_0;
  wire [1:0] simp4551_0;
  wire [1:0] simp4561_0;
  wire [7:0] fa3_25min_0;
  wire [1:0] simp4681_0;
  wire [1:0] simp4691_0;
  wire [7:0] fa3_26min_0;
  wire [1:0] simp4811_0;
  wire [1:0] simp4821_0;
  wire [7:0] fa3_27min_0;
  wire [1:0] simp4941_0;
  wire [1:0] simp4951_0;
  wire [7:0] fa3_28min_0;
  wire [1:0] simp5071_0;
  wire [1:0] simp5081_0;
  wire [7:0] fa3_29min_0;
  wire [1:0] simp5201_0;
  wire [1:0] simp5211_0;
  wire [7:0] fa3_30min_0;
  wire [1:0] simp5331_0;
  wire [1:0] simp5341_0;
  wire [7:0] fa3_31min_0;
  wire [1:0] simp5461_0;
  wire [1:0] simp5471_0;
  wire [7:0] fa3_32min_0;
  wire [1:0] simp5591_0;
  wire [1:0] simp5601_0;
  BUFF I0 (termf_1[0:0], i_0r0[0:0]);
  BUFF I1 (termf_1[1:1], i_0r0[1:1]);
  BUFF I2 (termf_1[2:2], i_0r0[2:2]);
  BUFF I3 (termf_1[3:3], i_0r0[3:3]);
  BUFF I4 (termf_1[4:4], i_0r0[4:4]);
  BUFF I5 (termf_1[5:5], i_0r0[5:5]);
  BUFF I6 (termf_1[6:6], i_0r0[6:6]);
  BUFF I7 (termf_1[7:7], i_0r0[7:7]);
  BUFF I8 (termf_1[8:8], i_0r0[8:8]);
  BUFF I9 (termf_1[9:9], i_0r0[9:9]);
  BUFF I10 (termf_1[10:10], i_0r0[10:10]);
  BUFF I11 (termf_1[11:11], i_0r0[11:11]);
  BUFF I12 (termf_1[12:12], i_0r0[12:12]);
  BUFF I13 (termf_1[13:13], i_0r0[13:13]);
  BUFF I14 (termf_1[14:14], i_0r0[14:14]);
  BUFF I15 (termf_1[15:15], i_0r0[15:15]);
  BUFF I16 (termf_1[16:16], i_0r0[16:16]);
  BUFF I17 (termf_1[17:17], i_0r0[17:17]);
  BUFF I18 (termf_1[18:18], i_0r0[18:18]);
  BUFF I19 (termf_1[19:19], i_0r0[19:19]);
  BUFF I20 (termf_1[20:20], i_0r0[20:20]);
  BUFF I21 (termf_1[21:21], i_0r0[21:21]);
  BUFF I22 (termf_1[22:22], i_0r0[22:22]);
  BUFF I23 (termf_1[23:23], i_0r0[23:23]);
  BUFF I24 (termf_1[24:24], i_0r0[24:24]);
  BUFF I25 (termf_1[25:25], i_0r0[25:25]);
  BUFF I26 (termf_1[26:26], i_0r0[26:26]);
  BUFF I27 (termf_1[27:27], i_0r0[27:27]);
  BUFF I28 (termf_1[28:28], i_0r0[28:28]);
  BUFF I29 (termf_1[29:29], i_0r0[29:29]);
  BUFF I30 (termf_1[30:30], i_0r0[30:30]);
  BUFF I31 (termf_1[31:31], i_0r0[31:31]);
  BUFF I32 (termf_1[32:32], i_0r0[31:31]);
  BUFF I33 (termt_1[0:0], i_0r1[0:0]);
  BUFF I34 (termt_1[1:1], i_0r1[1:1]);
  BUFF I35 (termt_1[2:2], i_0r1[2:2]);
  BUFF I36 (termt_1[3:3], i_0r1[3:3]);
  BUFF I37 (termt_1[4:4], i_0r1[4:4]);
  BUFF I38 (termt_1[5:5], i_0r1[5:5]);
  BUFF I39 (termt_1[6:6], i_0r1[6:6]);
  BUFF I40 (termt_1[7:7], i_0r1[7:7]);
  BUFF I41 (termt_1[8:8], i_0r1[8:8]);
  BUFF I42 (termt_1[9:9], i_0r1[9:9]);
  BUFF I43 (termt_1[10:10], i_0r1[10:10]);
  BUFF I44 (termt_1[11:11], i_0r1[11:11]);
  BUFF I45 (termt_1[12:12], i_0r1[12:12]);
  BUFF I46 (termt_1[13:13], i_0r1[13:13]);
  BUFF I47 (termt_1[14:14], i_0r1[14:14]);
  BUFF I48 (termt_1[15:15], i_0r1[15:15]);
  BUFF I49 (termt_1[16:16], i_0r1[16:16]);
  BUFF I50 (termt_1[17:17], i_0r1[17:17]);
  BUFF I51 (termt_1[18:18], i_0r1[18:18]);
  BUFF I52 (termt_1[19:19], i_0r1[19:19]);
  BUFF I53 (termt_1[20:20], i_0r1[20:20]);
  BUFF I54 (termt_1[21:21], i_0r1[21:21]);
  BUFF I55 (termt_1[22:22], i_0r1[22:22]);
  BUFF I56 (termt_1[23:23], i_0r1[23:23]);
  BUFF I57 (termt_1[24:24], i_0r1[24:24]);
  BUFF I58 (termt_1[25:25], i_0r1[25:25]);
  BUFF I59 (termt_1[26:26], i_0r1[26:26]);
  BUFF I60 (termt_1[27:27], i_0r1[27:27]);
  BUFF I61 (termt_1[28:28], i_0r1[28:28]);
  BUFF I62 (termt_1[29:29], i_0r1[29:29]);
  BUFF I63 (termt_1[30:30], i_0r1[30:30]);
  BUFF I64 (termt_1[31:31], i_0r1[31:31]);
  BUFF I65 (termt_1[32:32], i_0r1[31:31]);
  BUFF I66 (termf_2[0:0], i_0r0[32:32]);
  BUFF I67 (termf_2[1:1], i_0r0[33:33]);
  BUFF I68 (termf_2[2:2], i_0r0[34:34]);
  BUFF I69 (termf_2[3:3], i_0r0[35:35]);
  BUFF I70 (termf_2[4:4], i_0r0[36:36]);
  BUFF I71 (termf_2[5:5], i_0r0[37:37]);
  BUFF I72 (termf_2[6:6], i_0r0[38:38]);
  BUFF I73 (termf_2[7:7], i_0r0[39:39]);
  BUFF I74 (termf_2[8:8], i_0r0[40:40]);
  BUFF I75 (termf_2[9:9], i_0r0[41:41]);
  BUFF I76 (termf_2[10:10], i_0r0[42:42]);
  BUFF I77 (termf_2[11:11], i_0r0[43:43]);
  BUFF I78 (termf_2[12:12], i_0r0[44:44]);
  BUFF I79 (termf_2[13:13], i_0r0[45:45]);
  BUFF I80 (termf_2[14:14], i_0r0[46:46]);
  BUFF I81 (termf_2[15:15], i_0r0[47:47]);
  BUFF I82 (termf_2[16:16], i_0r0[48:48]);
  BUFF I83 (termf_2[17:17], i_0r0[49:49]);
  BUFF I84 (termf_2[18:18], i_0r0[50:50]);
  BUFF I85 (termf_2[19:19], i_0r0[51:51]);
  BUFF I86 (termf_2[20:20], i_0r0[52:52]);
  BUFF I87 (termf_2[21:21], i_0r0[53:53]);
  BUFF I88 (termf_2[22:22], i_0r0[54:54]);
  BUFF I89 (termf_2[23:23], i_0r0[55:55]);
  BUFF I90 (termf_2[24:24], i_0r0[56:56]);
  BUFF I91 (termf_2[25:25], i_0r0[57:57]);
  BUFF I92 (termf_2[26:26], i_0r0[58:58]);
  BUFF I93 (termf_2[27:27], i_0r0[59:59]);
  BUFF I94 (termf_2[28:28], i_0r0[60:60]);
  BUFF I95 (termf_2[29:29], i_0r0[61:61]);
  BUFF I96 (termf_2[30:30], i_0r0[62:62]);
  BUFF I97 (termf_2[31:31], i_0r0[63:63]);
  BUFF I98 (termf_2[32:32], i_0r0[63:63]);
  BUFF I99 (termt_2[0:0], i_0r1[32:32]);
  BUFF I100 (termt_2[1:1], i_0r1[33:33]);
  BUFF I101 (termt_2[2:2], i_0r1[34:34]);
  BUFF I102 (termt_2[3:3], i_0r1[35:35]);
  BUFF I103 (termt_2[4:4], i_0r1[36:36]);
  BUFF I104 (termt_2[5:5], i_0r1[37:37]);
  BUFF I105 (termt_2[6:6], i_0r1[38:38]);
  BUFF I106 (termt_2[7:7], i_0r1[39:39]);
  BUFF I107 (termt_2[8:8], i_0r1[40:40]);
  BUFF I108 (termt_2[9:9], i_0r1[41:41]);
  BUFF I109 (termt_2[10:10], i_0r1[42:42]);
  BUFF I110 (termt_2[11:11], i_0r1[43:43]);
  BUFF I111 (termt_2[12:12], i_0r1[44:44]);
  BUFF I112 (termt_2[13:13], i_0r1[45:45]);
  BUFF I113 (termt_2[14:14], i_0r1[46:46]);
  BUFF I114 (termt_2[15:15], i_0r1[47:47]);
  BUFF I115 (termt_2[16:16], i_0r1[48:48]);
  BUFF I116 (termt_2[17:17], i_0r1[49:49]);
  BUFF I117 (termt_2[18:18], i_0r1[50:50]);
  BUFF I118 (termt_2[19:19], i_0r1[51:51]);
  BUFF I119 (termt_2[20:20], i_0r1[52:52]);
  BUFF I120 (termt_2[21:21], i_0r1[53:53]);
  BUFF I121 (termt_2[22:22], i_0r1[54:54]);
  BUFF I122 (termt_2[23:23], i_0r1[55:55]);
  BUFF I123 (termt_2[24:24], i_0r1[56:56]);
  BUFF I124 (termt_2[25:25], i_0r1[57:57]);
  BUFF I125 (termt_2[26:26], i_0r1[58:58]);
  BUFF I126 (termt_2[27:27], i_0r1[59:59]);
  BUFF I127 (termt_2[28:28], i_0r1[60:60]);
  BUFF I128 (termt_2[29:29], i_0r1[61:61]);
  BUFF I129 (termt_2[30:30], i_0r1[62:62]);
  BUFF I130 (termt_2[31:31], i_0r1[63:63]);
  BUFF I131 (termt_2[32:32], i_0r1[63:63]);
  C2 I132 (ha3__0[0:0], termf_2[0:0], termf_1[0:0]);
  C2 I133 (ha3__0[1:1], termf_2[0:0], termt_1[0:0]);
  C2 I134 (ha3__0[2:2], termt_2[0:0], termf_1[0:0]);
  C2 I135 (ha3__0[3:3], termt_2[0:0], termt_1[0:0]);
  OR3 I136 (cf3__0[0:0], ha3__0[0:0], ha3__0[1:1], ha3__0[2:2]);
  BUFF I137 (ct3__0[0:0], ha3__0[3:3]);
  OR2 I138 (o_0r0[0:0], ha3__0[0:0], ha3__0[3:3]);
  OR2 I139 (o_0r1[0:0], ha3__0[1:1], ha3__0[2:2]);
  C3 I140 (fa3_1min_0[0:0], cf3__0[0:0], termf_2[1:1], termf_1[1:1]);
  C3 I141 (fa3_1min_0[1:1], cf3__0[0:0], termf_2[1:1], termt_1[1:1]);
  C3 I142 (fa3_1min_0[2:2], cf3__0[0:0], termt_2[1:1], termf_1[1:1]);
  C3 I143 (fa3_1min_0[3:3], cf3__0[0:0], termt_2[1:1], termt_1[1:1]);
  C3 I144 (fa3_1min_0[4:4], ct3__0[0:0], termf_2[1:1], termf_1[1:1]);
  C3 I145 (fa3_1min_0[5:5], ct3__0[0:0], termf_2[1:1], termt_1[1:1]);
  C3 I146 (fa3_1min_0[6:6], ct3__0[0:0], termt_2[1:1], termf_1[1:1]);
  C3 I147 (fa3_1min_0[7:7], ct3__0[0:0], termt_2[1:1], termt_1[1:1]);
  NOR3 I148 (simp1561_0[0:0], fa3_1min_0[0:0], fa3_1min_0[3:3], fa3_1min_0[5:5]);
  INV I149 (simp1561_0[1:1], fa3_1min_0[6:6]);
  NAND2 I150 (o_0r0[1:1], simp1561_0[0:0], simp1561_0[1:1]);
  NOR3 I151 (simp1571_0[0:0], fa3_1min_0[1:1], fa3_1min_0[2:2], fa3_1min_0[4:4]);
  INV I152 (simp1571_0[1:1], fa3_1min_0[7:7]);
  NAND2 I153 (o_0r1[1:1], simp1571_0[0:0], simp1571_0[1:1]);
  AO222 I154 (ct3__0[1:1], termt_1[1:1], termt_2[1:1], termt_1[1:1], ct3__0[0:0], termt_2[1:1], ct3__0[0:0]);
  AO222 I155 (cf3__0[1:1], termf_1[1:1], termf_2[1:1], termf_1[1:1], cf3__0[0:0], termf_2[1:1], cf3__0[0:0]);
  C3 I156 (fa3_2min_0[0:0], cf3__0[1:1], termf_2[2:2], termf_1[2:2]);
  C3 I157 (fa3_2min_0[1:1], cf3__0[1:1], termf_2[2:2], termt_1[2:2]);
  C3 I158 (fa3_2min_0[2:2], cf3__0[1:1], termt_2[2:2], termf_1[2:2]);
  C3 I159 (fa3_2min_0[3:3], cf3__0[1:1], termt_2[2:2], termt_1[2:2]);
  C3 I160 (fa3_2min_0[4:4], ct3__0[1:1], termf_2[2:2], termf_1[2:2]);
  C3 I161 (fa3_2min_0[5:5], ct3__0[1:1], termf_2[2:2], termt_1[2:2]);
  C3 I162 (fa3_2min_0[6:6], ct3__0[1:1], termt_2[2:2], termf_1[2:2]);
  C3 I163 (fa3_2min_0[7:7], ct3__0[1:1], termt_2[2:2], termt_1[2:2]);
  NOR3 I164 (simp1691_0[0:0], fa3_2min_0[0:0], fa3_2min_0[3:3], fa3_2min_0[5:5]);
  INV I165 (simp1691_0[1:1], fa3_2min_0[6:6]);
  NAND2 I166 (o_0r0[2:2], simp1691_0[0:0], simp1691_0[1:1]);
  NOR3 I167 (simp1701_0[0:0], fa3_2min_0[1:1], fa3_2min_0[2:2], fa3_2min_0[4:4]);
  INV I168 (simp1701_0[1:1], fa3_2min_0[7:7]);
  NAND2 I169 (o_0r1[2:2], simp1701_0[0:0], simp1701_0[1:1]);
  AO222 I170 (ct3__0[2:2], termt_1[2:2], termt_2[2:2], termt_1[2:2], ct3__0[1:1], termt_2[2:2], ct3__0[1:1]);
  AO222 I171 (cf3__0[2:2], termf_1[2:2], termf_2[2:2], termf_1[2:2], cf3__0[1:1], termf_2[2:2], cf3__0[1:1]);
  C3 I172 (fa3_3min_0[0:0], cf3__0[2:2], termf_2[3:3], termf_1[3:3]);
  C3 I173 (fa3_3min_0[1:1], cf3__0[2:2], termf_2[3:3], termt_1[3:3]);
  C3 I174 (fa3_3min_0[2:2], cf3__0[2:2], termt_2[3:3], termf_1[3:3]);
  C3 I175 (fa3_3min_0[3:3], cf3__0[2:2], termt_2[3:3], termt_1[3:3]);
  C3 I176 (fa3_3min_0[4:4], ct3__0[2:2], termf_2[3:3], termf_1[3:3]);
  C3 I177 (fa3_3min_0[5:5], ct3__0[2:2], termf_2[3:3], termt_1[3:3]);
  C3 I178 (fa3_3min_0[6:6], ct3__0[2:2], termt_2[3:3], termf_1[3:3]);
  C3 I179 (fa3_3min_0[7:7], ct3__0[2:2], termt_2[3:3], termt_1[3:3]);
  NOR3 I180 (simp1821_0[0:0], fa3_3min_0[0:0], fa3_3min_0[3:3], fa3_3min_0[5:5]);
  INV I181 (simp1821_0[1:1], fa3_3min_0[6:6]);
  NAND2 I182 (o_0r0[3:3], simp1821_0[0:0], simp1821_0[1:1]);
  NOR3 I183 (simp1831_0[0:0], fa3_3min_0[1:1], fa3_3min_0[2:2], fa3_3min_0[4:4]);
  INV I184 (simp1831_0[1:1], fa3_3min_0[7:7]);
  NAND2 I185 (o_0r1[3:3], simp1831_0[0:0], simp1831_0[1:1]);
  AO222 I186 (ct3__0[3:3], termt_1[3:3], termt_2[3:3], termt_1[3:3], ct3__0[2:2], termt_2[3:3], ct3__0[2:2]);
  AO222 I187 (cf3__0[3:3], termf_1[3:3], termf_2[3:3], termf_1[3:3], cf3__0[2:2], termf_2[3:3], cf3__0[2:2]);
  C3 I188 (fa3_4min_0[0:0], cf3__0[3:3], termf_2[4:4], termf_1[4:4]);
  C3 I189 (fa3_4min_0[1:1], cf3__0[3:3], termf_2[4:4], termt_1[4:4]);
  C3 I190 (fa3_4min_0[2:2], cf3__0[3:3], termt_2[4:4], termf_1[4:4]);
  C3 I191 (fa3_4min_0[3:3], cf3__0[3:3], termt_2[4:4], termt_1[4:4]);
  C3 I192 (fa3_4min_0[4:4], ct3__0[3:3], termf_2[4:4], termf_1[4:4]);
  C3 I193 (fa3_4min_0[5:5], ct3__0[3:3], termf_2[4:4], termt_1[4:4]);
  C3 I194 (fa3_4min_0[6:6], ct3__0[3:3], termt_2[4:4], termf_1[4:4]);
  C3 I195 (fa3_4min_0[7:7], ct3__0[3:3], termt_2[4:4], termt_1[4:4]);
  NOR3 I196 (simp1951_0[0:0], fa3_4min_0[0:0], fa3_4min_0[3:3], fa3_4min_0[5:5]);
  INV I197 (simp1951_0[1:1], fa3_4min_0[6:6]);
  NAND2 I198 (o_0r0[4:4], simp1951_0[0:0], simp1951_0[1:1]);
  NOR3 I199 (simp1961_0[0:0], fa3_4min_0[1:1], fa3_4min_0[2:2], fa3_4min_0[4:4]);
  INV I200 (simp1961_0[1:1], fa3_4min_0[7:7]);
  NAND2 I201 (o_0r1[4:4], simp1961_0[0:0], simp1961_0[1:1]);
  AO222 I202 (ct3__0[4:4], termt_1[4:4], termt_2[4:4], termt_1[4:4], ct3__0[3:3], termt_2[4:4], ct3__0[3:3]);
  AO222 I203 (cf3__0[4:4], termf_1[4:4], termf_2[4:4], termf_1[4:4], cf3__0[3:3], termf_2[4:4], cf3__0[3:3]);
  C3 I204 (fa3_5min_0[0:0], cf3__0[4:4], termf_2[5:5], termf_1[5:5]);
  C3 I205 (fa3_5min_0[1:1], cf3__0[4:4], termf_2[5:5], termt_1[5:5]);
  C3 I206 (fa3_5min_0[2:2], cf3__0[4:4], termt_2[5:5], termf_1[5:5]);
  C3 I207 (fa3_5min_0[3:3], cf3__0[4:4], termt_2[5:5], termt_1[5:5]);
  C3 I208 (fa3_5min_0[4:4], ct3__0[4:4], termf_2[5:5], termf_1[5:5]);
  C3 I209 (fa3_5min_0[5:5], ct3__0[4:4], termf_2[5:5], termt_1[5:5]);
  C3 I210 (fa3_5min_0[6:6], ct3__0[4:4], termt_2[5:5], termf_1[5:5]);
  C3 I211 (fa3_5min_0[7:7], ct3__0[4:4], termt_2[5:5], termt_1[5:5]);
  NOR3 I212 (simp2081_0[0:0], fa3_5min_0[0:0], fa3_5min_0[3:3], fa3_5min_0[5:5]);
  INV I213 (simp2081_0[1:1], fa3_5min_0[6:6]);
  NAND2 I214 (o_0r0[5:5], simp2081_0[0:0], simp2081_0[1:1]);
  NOR3 I215 (simp2091_0[0:0], fa3_5min_0[1:1], fa3_5min_0[2:2], fa3_5min_0[4:4]);
  INV I216 (simp2091_0[1:1], fa3_5min_0[7:7]);
  NAND2 I217 (o_0r1[5:5], simp2091_0[0:0], simp2091_0[1:1]);
  AO222 I218 (ct3__0[5:5], termt_1[5:5], termt_2[5:5], termt_1[5:5], ct3__0[4:4], termt_2[5:5], ct3__0[4:4]);
  AO222 I219 (cf3__0[5:5], termf_1[5:5], termf_2[5:5], termf_1[5:5], cf3__0[4:4], termf_2[5:5], cf3__0[4:4]);
  C3 I220 (fa3_6min_0[0:0], cf3__0[5:5], termf_2[6:6], termf_1[6:6]);
  C3 I221 (fa3_6min_0[1:1], cf3__0[5:5], termf_2[6:6], termt_1[6:6]);
  C3 I222 (fa3_6min_0[2:2], cf3__0[5:5], termt_2[6:6], termf_1[6:6]);
  C3 I223 (fa3_6min_0[3:3], cf3__0[5:5], termt_2[6:6], termt_1[6:6]);
  C3 I224 (fa3_6min_0[4:4], ct3__0[5:5], termf_2[6:6], termf_1[6:6]);
  C3 I225 (fa3_6min_0[5:5], ct3__0[5:5], termf_2[6:6], termt_1[6:6]);
  C3 I226 (fa3_6min_0[6:6], ct3__0[5:5], termt_2[6:6], termf_1[6:6]);
  C3 I227 (fa3_6min_0[7:7], ct3__0[5:5], termt_2[6:6], termt_1[6:6]);
  NOR3 I228 (simp2211_0[0:0], fa3_6min_0[0:0], fa3_6min_0[3:3], fa3_6min_0[5:5]);
  INV I229 (simp2211_0[1:1], fa3_6min_0[6:6]);
  NAND2 I230 (o_0r0[6:6], simp2211_0[0:0], simp2211_0[1:1]);
  NOR3 I231 (simp2221_0[0:0], fa3_6min_0[1:1], fa3_6min_0[2:2], fa3_6min_0[4:4]);
  INV I232 (simp2221_0[1:1], fa3_6min_0[7:7]);
  NAND2 I233 (o_0r1[6:6], simp2221_0[0:0], simp2221_0[1:1]);
  AO222 I234 (ct3__0[6:6], termt_1[6:6], termt_2[6:6], termt_1[6:6], ct3__0[5:5], termt_2[6:6], ct3__0[5:5]);
  AO222 I235 (cf3__0[6:6], termf_1[6:6], termf_2[6:6], termf_1[6:6], cf3__0[5:5], termf_2[6:6], cf3__0[5:5]);
  C3 I236 (fa3_7min_0[0:0], cf3__0[6:6], termf_2[7:7], termf_1[7:7]);
  C3 I237 (fa3_7min_0[1:1], cf3__0[6:6], termf_2[7:7], termt_1[7:7]);
  C3 I238 (fa3_7min_0[2:2], cf3__0[6:6], termt_2[7:7], termf_1[7:7]);
  C3 I239 (fa3_7min_0[3:3], cf3__0[6:6], termt_2[7:7], termt_1[7:7]);
  C3 I240 (fa3_7min_0[4:4], ct3__0[6:6], termf_2[7:7], termf_1[7:7]);
  C3 I241 (fa3_7min_0[5:5], ct3__0[6:6], termf_2[7:7], termt_1[7:7]);
  C3 I242 (fa3_7min_0[6:6], ct3__0[6:6], termt_2[7:7], termf_1[7:7]);
  C3 I243 (fa3_7min_0[7:7], ct3__0[6:6], termt_2[7:7], termt_1[7:7]);
  NOR3 I244 (simp2341_0[0:0], fa3_7min_0[0:0], fa3_7min_0[3:3], fa3_7min_0[5:5]);
  INV I245 (simp2341_0[1:1], fa3_7min_0[6:6]);
  NAND2 I246 (o_0r0[7:7], simp2341_0[0:0], simp2341_0[1:1]);
  NOR3 I247 (simp2351_0[0:0], fa3_7min_0[1:1], fa3_7min_0[2:2], fa3_7min_0[4:4]);
  INV I248 (simp2351_0[1:1], fa3_7min_0[7:7]);
  NAND2 I249 (o_0r1[7:7], simp2351_0[0:0], simp2351_0[1:1]);
  AO222 I250 (ct3__0[7:7], termt_1[7:7], termt_2[7:7], termt_1[7:7], ct3__0[6:6], termt_2[7:7], ct3__0[6:6]);
  AO222 I251 (cf3__0[7:7], termf_1[7:7], termf_2[7:7], termf_1[7:7], cf3__0[6:6], termf_2[7:7], cf3__0[6:6]);
  C3 I252 (fa3_8min_0[0:0], cf3__0[7:7], termf_2[8:8], termf_1[8:8]);
  C3 I253 (fa3_8min_0[1:1], cf3__0[7:7], termf_2[8:8], termt_1[8:8]);
  C3 I254 (fa3_8min_0[2:2], cf3__0[7:7], termt_2[8:8], termf_1[8:8]);
  C3 I255 (fa3_8min_0[3:3], cf3__0[7:7], termt_2[8:8], termt_1[8:8]);
  C3 I256 (fa3_8min_0[4:4], ct3__0[7:7], termf_2[8:8], termf_1[8:8]);
  C3 I257 (fa3_8min_0[5:5], ct3__0[7:7], termf_2[8:8], termt_1[8:8]);
  C3 I258 (fa3_8min_0[6:6], ct3__0[7:7], termt_2[8:8], termf_1[8:8]);
  C3 I259 (fa3_8min_0[7:7], ct3__0[7:7], termt_2[8:8], termt_1[8:8]);
  NOR3 I260 (simp2471_0[0:0], fa3_8min_0[0:0], fa3_8min_0[3:3], fa3_8min_0[5:5]);
  INV I261 (simp2471_0[1:1], fa3_8min_0[6:6]);
  NAND2 I262 (o_0r0[8:8], simp2471_0[0:0], simp2471_0[1:1]);
  NOR3 I263 (simp2481_0[0:0], fa3_8min_0[1:1], fa3_8min_0[2:2], fa3_8min_0[4:4]);
  INV I264 (simp2481_0[1:1], fa3_8min_0[7:7]);
  NAND2 I265 (o_0r1[8:8], simp2481_0[0:0], simp2481_0[1:1]);
  AO222 I266 (ct3__0[8:8], termt_1[8:8], termt_2[8:8], termt_1[8:8], ct3__0[7:7], termt_2[8:8], ct3__0[7:7]);
  AO222 I267 (cf3__0[8:8], termf_1[8:8], termf_2[8:8], termf_1[8:8], cf3__0[7:7], termf_2[8:8], cf3__0[7:7]);
  C3 I268 (fa3_9min_0[0:0], cf3__0[8:8], termf_2[9:9], termf_1[9:9]);
  C3 I269 (fa3_9min_0[1:1], cf3__0[8:8], termf_2[9:9], termt_1[9:9]);
  C3 I270 (fa3_9min_0[2:2], cf3__0[8:8], termt_2[9:9], termf_1[9:9]);
  C3 I271 (fa3_9min_0[3:3], cf3__0[8:8], termt_2[9:9], termt_1[9:9]);
  C3 I272 (fa3_9min_0[4:4], ct3__0[8:8], termf_2[9:9], termf_1[9:9]);
  C3 I273 (fa3_9min_0[5:5], ct3__0[8:8], termf_2[9:9], termt_1[9:9]);
  C3 I274 (fa3_9min_0[6:6], ct3__0[8:8], termt_2[9:9], termf_1[9:9]);
  C3 I275 (fa3_9min_0[7:7], ct3__0[8:8], termt_2[9:9], termt_1[9:9]);
  NOR3 I276 (simp2601_0[0:0], fa3_9min_0[0:0], fa3_9min_0[3:3], fa3_9min_0[5:5]);
  INV I277 (simp2601_0[1:1], fa3_9min_0[6:6]);
  NAND2 I278 (o_0r0[9:9], simp2601_0[0:0], simp2601_0[1:1]);
  NOR3 I279 (simp2611_0[0:0], fa3_9min_0[1:1], fa3_9min_0[2:2], fa3_9min_0[4:4]);
  INV I280 (simp2611_0[1:1], fa3_9min_0[7:7]);
  NAND2 I281 (o_0r1[9:9], simp2611_0[0:0], simp2611_0[1:1]);
  AO222 I282 (ct3__0[9:9], termt_1[9:9], termt_2[9:9], termt_1[9:9], ct3__0[8:8], termt_2[9:9], ct3__0[8:8]);
  AO222 I283 (cf3__0[9:9], termf_1[9:9], termf_2[9:9], termf_1[9:9], cf3__0[8:8], termf_2[9:9], cf3__0[8:8]);
  C3 I284 (fa3_10min_0[0:0], cf3__0[9:9], termf_2[10:10], termf_1[10:10]);
  C3 I285 (fa3_10min_0[1:1], cf3__0[9:9], termf_2[10:10], termt_1[10:10]);
  C3 I286 (fa3_10min_0[2:2], cf3__0[9:9], termt_2[10:10], termf_1[10:10]);
  C3 I287 (fa3_10min_0[3:3], cf3__0[9:9], termt_2[10:10], termt_1[10:10]);
  C3 I288 (fa3_10min_0[4:4], ct3__0[9:9], termf_2[10:10], termf_1[10:10]);
  C3 I289 (fa3_10min_0[5:5], ct3__0[9:9], termf_2[10:10], termt_1[10:10]);
  C3 I290 (fa3_10min_0[6:6], ct3__0[9:9], termt_2[10:10], termf_1[10:10]);
  C3 I291 (fa3_10min_0[7:7], ct3__0[9:9], termt_2[10:10], termt_1[10:10]);
  NOR3 I292 (simp2731_0[0:0], fa3_10min_0[0:0], fa3_10min_0[3:3], fa3_10min_0[5:5]);
  INV I293 (simp2731_0[1:1], fa3_10min_0[6:6]);
  NAND2 I294 (o_0r0[10:10], simp2731_0[0:0], simp2731_0[1:1]);
  NOR3 I295 (simp2741_0[0:0], fa3_10min_0[1:1], fa3_10min_0[2:2], fa3_10min_0[4:4]);
  INV I296 (simp2741_0[1:1], fa3_10min_0[7:7]);
  NAND2 I297 (o_0r1[10:10], simp2741_0[0:0], simp2741_0[1:1]);
  AO222 I298 (ct3__0[10:10], termt_1[10:10], termt_2[10:10], termt_1[10:10], ct3__0[9:9], termt_2[10:10], ct3__0[9:9]);
  AO222 I299 (cf3__0[10:10], termf_1[10:10], termf_2[10:10], termf_1[10:10], cf3__0[9:9], termf_2[10:10], cf3__0[9:9]);
  C3 I300 (fa3_11min_0[0:0], cf3__0[10:10], termf_2[11:11], termf_1[11:11]);
  C3 I301 (fa3_11min_0[1:1], cf3__0[10:10], termf_2[11:11], termt_1[11:11]);
  C3 I302 (fa3_11min_0[2:2], cf3__0[10:10], termt_2[11:11], termf_1[11:11]);
  C3 I303 (fa3_11min_0[3:3], cf3__0[10:10], termt_2[11:11], termt_1[11:11]);
  C3 I304 (fa3_11min_0[4:4], ct3__0[10:10], termf_2[11:11], termf_1[11:11]);
  C3 I305 (fa3_11min_0[5:5], ct3__0[10:10], termf_2[11:11], termt_1[11:11]);
  C3 I306 (fa3_11min_0[6:6], ct3__0[10:10], termt_2[11:11], termf_1[11:11]);
  C3 I307 (fa3_11min_0[7:7], ct3__0[10:10], termt_2[11:11], termt_1[11:11]);
  NOR3 I308 (simp2861_0[0:0], fa3_11min_0[0:0], fa3_11min_0[3:3], fa3_11min_0[5:5]);
  INV I309 (simp2861_0[1:1], fa3_11min_0[6:6]);
  NAND2 I310 (o_0r0[11:11], simp2861_0[0:0], simp2861_0[1:1]);
  NOR3 I311 (simp2871_0[0:0], fa3_11min_0[1:1], fa3_11min_0[2:2], fa3_11min_0[4:4]);
  INV I312 (simp2871_0[1:1], fa3_11min_0[7:7]);
  NAND2 I313 (o_0r1[11:11], simp2871_0[0:0], simp2871_0[1:1]);
  AO222 I314 (ct3__0[11:11], termt_1[11:11], termt_2[11:11], termt_1[11:11], ct3__0[10:10], termt_2[11:11], ct3__0[10:10]);
  AO222 I315 (cf3__0[11:11], termf_1[11:11], termf_2[11:11], termf_1[11:11], cf3__0[10:10], termf_2[11:11], cf3__0[10:10]);
  C3 I316 (fa3_12min_0[0:0], cf3__0[11:11], termf_2[12:12], termf_1[12:12]);
  C3 I317 (fa3_12min_0[1:1], cf3__0[11:11], termf_2[12:12], termt_1[12:12]);
  C3 I318 (fa3_12min_0[2:2], cf3__0[11:11], termt_2[12:12], termf_1[12:12]);
  C3 I319 (fa3_12min_0[3:3], cf3__0[11:11], termt_2[12:12], termt_1[12:12]);
  C3 I320 (fa3_12min_0[4:4], ct3__0[11:11], termf_2[12:12], termf_1[12:12]);
  C3 I321 (fa3_12min_0[5:5], ct3__0[11:11], termf_2[12:12], termt_1[12:12]);
  C3 I322 (fa3_12min_0[6:6], ct3__0[11:11], termt_2[12:12], termf_1[12:12]);
  C3 I323 (fa3_12min_0[7:7], ct3__0[11:11], termt_2[12:12], termt_1[12:12]);
  NOR3 I324 (simp2991_0[0:0], fa3_12min_0[0:0], fa3_12min_0[3:3], fa3_12min_0[5:5]);
  INV I325 (simp2991_0[1:1], fa3_12min_0[6:6]);
  NAND2 I326 (o_0r0[12:12], simp2991_0[0:0], simp2991_0[1:1]);
  NOR3 I327 (simp3001_0[0:0], fa3_12min_0[1:1], fa3_12min_0[2:2], fa3_12min_0[4:4]);
  INV I328 (simp3001_0[1:1], fa3_12min_0[7:7]);
  NAND2 I329 (o_0r1[12:12], simp3001_0[0:0], simp3001_0[1:1]);
  AO222 I330 (ct3__0[12:12], termt_1[12:12], termt_2[12:12], termt_1[12:12], ct3__0[11:11], termt_2[12:12], ct3__0[11:11]);
  AO222 I331 (cf3__0[12:12], termf_1[12:12], termf_2[12:12], termf_1[12:12], cf3__0[11:11], termf_2[12:12], cf3__0[11:11]);
  C3 I332 (fa3_13min_0[0:0], cf3__0[12:12], termf_2[13:13], termf_1[13:13]);
  C3 I333 (fa3_13min_0[1:1], cf3__0[12:12], termf_2[13:13], termt_1[13:13]);
  C3 I334 (fa3_13min_0[2:2], cf3__0[12:12], termt_2[13:13], termf_1[13:13]);
  C3 I335 (fa3_13min_0[3:3], cf3__0[12:12], termt_2[13:13], termt_1[13:13]);
  C3 I336 (fa3_13min_0[4:4], ct3__0[12:12], termf_2[13:13], termf_1[13:13]);
  C3 I337 (fa3_13min_0[5:5], ct3__0[12:12], termf_2[13:13], termt_1[13:13]);
  C3 I338 (fa3_13min_0[6:6], ct3__0[12:12], termt_2[13:13], termf_1[13:13]);
  C3 I339 (fa3_13min_0[7:7], ct3__0[12:12], termt_2[13:13], termt_1[13:13]);
  NOR3 I340 (simp3121_0[0:0], fa3_13min_0[0:0], fa3_13min_0[3:3], fa3_13min_0[5:5]);
  INV I341 (simp3121_0[1:1], fa3_13min_0[6:6]);
  NAND2 I342 (o_0r0[13:13], simp3121_0[0:0], simp3121_0[1:1]);
  NOR3 I343 (simp3131_0[0:0], fa3_13min_0[1:1], fa3_13min_0[2:2], fa3_13min_0[4:4]);
  INV I344 (simp3131_0[1:1], fa3_13min_0[7:7]);
  NAND2 I345 (o_0r1[13:13], simp3131_0[0:0], simp3131_0[1:1]);
  AO222 I346 (ct3__0[13:13], termt_1[13:13], termt_2[13:13], termt_1[13:13], ct3__0[12:12], termt_2[13:13], ct3__0[12:12]);
  AO222 I347 (cf3__0[13:13], termf_1[13:13], termf_2[13:13], termf_1[13:13], cf3__0[12:12], termf_2[13:13], cf3__0[12:12]);
  C3 I348 (fa3_14min_0[0:0], cf3__0[13:13], termf_2[14:14], termf_1[14:14]);
  C3 I349 (fa3_14min_0[1:1], cf3__0[13:13], termf_2[14:14], termt_1[14:14]);
  C3 I350 (fa3_14min_0[2:2], cf3__0[13:13], termt_2[14:14], termf_1[14:14]);
  C3 I351 (fa3_14min_0[3:3], cf3__0[13:13], termt_2[14:14], termt_1[14:14]);
  C3 I352 (fa3_14min_0[4:4], ct3__0[13:13], termf_2[14:14], termf_1[14:14]);
  C3 I353 (fa3_14min_0[5:5], ct3__0[13:13], termf_2[14:14], termt_1[14:14]);
  C3 I354 (fa3_14min_0[6:6], ct3__0[13:13], termt_2[14:14], termf_1[14:14]);
  C3 I355 (fa3_14min_0[7:7], ct3__0[13:13], termt_2[14:14], termt_1[14:14]);
  NOR3 I356 (simp3251_0[0:0], fa3_14min_0[0:0], fa3_14min_0[3:3], fa3_14min_0[5:5]);
  INV I357 (simp3251_0[1:1], fa3_14min_0[6:6]);
  NAND2 I358 (o_0r0[14:14], simp3251_0[0:0], simp3251_0[1:1]);
  NOR3 I359 (simp3261_0[0:0], fa3_14min_0[1:1], fa3_14min_0[2:2], fa3_14min_0[4:4]);
  INV I360 (simp3261_0[1:1], fa3_14min_0[7:7]);
  NAND2 I361 (o_0r1[14:14], simp3261_0[0:0], simp3261_0[1:1]);
  AO222 I362 (ct3__0[14:14], termt_1[14:14], termt_2[14:14], termt_1[14:14], ct3__0[13:13], termt_2[14:14], ct3__0[13:13]);
  AO222 I363 (cf3__0[14:14], termf_1[14:14], termf_2[14:14], termf_1[14:14], cf3__0[13:13], termf_2[14:14], cf3__0[13:13]);
  C3 I364 (fa3_15min_0[0:0], cf3__0[14:14], termf_2[15:15], termf_1[15:15]);
  C3 I365 (fa3_15min_0[1:1], cf3__0[14:14], termf_2[15:15], termt_1[15:15]);
  C3 I366 (fa3_15min_0[2:2], cf3__0[14:14], termt_2[15:15], termf_1[15:15]);
  C3 I367 (fa3_15min_0[3:3], cf3__0[14:14], termt_2[15:15], termt_1[15:15]);
  C3 I368 (fa3_15min_0[4:4], ct3__0[14:14], termf_2[15:15], termf_1[15:15]);
  C3 I369 (fa3_15min_0[5:5], ct3__0[14:14], termf_2[15:15], termt_1[15:15]);
  C3 I370 (fa3_15min_0[6:6], ct3__0[14:14], termt_2[15:15], termf_1[15:15]);
  C3 I371 (fa3_15min_0[7:7], ct3__0[14:14], termt_2[15:15], termt_1[15:15]);
  NOR3 I372 (simp3381_0[0:0], fa3_15min_0[0:0], fa3_15min_0[3:3], fa3_15min_0[5:5]);
  INV I373 (simp3381_0[1:1], fa3_15min_0[6:6]);
  NAND2 I374 (o_0r0[15:15], simp3381_0[0:0], simp3381_0[1:1]);
  NOR3 I375 (simp3391_0[0:0], fa3_15min_0[1:1], fa3_15min_0[2:2], fa3_15min_0[4:4]);
  INV I376 (simp3391_0[1:1], fa3_15min_0[7:7]);
  NAND2 I377 (o_0r1[15:15], simp3391_0[0:0], simp3391_0[1:1]);
  AO222 I378 (ct3__0[15:15], termt_1[15:15], termt_2[15:15], termt_1[15:15], ct3__0[14:14], termt_2[15:15], ct3__0[14:14]);
  AO222 I379 (cf3__0[15:15], termf_1[15:15], termf_2[15:15], termf_1[15:15], cf3__0[14:14], termf_2[15:15], cf3__0[14:14]);
  C3 I380 (fa3_16min_0[0:0], cf3__0[15:15], termf_2[16:16], termf_1[16:16]);
  C3 I381 (fa3_16min_0[1:1], cf3__0[15:15], termf_2[16:16], termt_1[16:16]);
  C3 I382 (fa3_16min_0[2:2], cf3__0[15:15], termt_2[16:16], termf_1[16:16]);
  C3 I383 (fa3_16min_0[3:3], cf3__0[15:15], termt_2[16:16], termt_1[16:16]);
  C3 I384 (fa3_16min_0[4:4], ct3__0[15:15], termf_2[16:16], termf_1[16:16]);
  C3 I385 (fa3_16min_0[5:5], ct3__0[15:15], termf_2[16:16], termt_1[16:16]);
  C3 I386 (fa3_16min_0[6:6], ct3__0[15:15], termt_2[16:16], termf_1[16:16]);
  C3 I387 (fa3_16min_0[7:7], ct3__0[15:15], termt_2[16:16], termt_1[16:16]);
  NOR3 I388 (simp3511_0[0:0], fa3_16min_0[0:0], fa3_16min_0[3:3], fa3_16min_0[5:5]);
  INV I389 (simp3511_0[1:1], fa3_16min_0[6:6]);
  NAND2 I390 (o_0r0[16:16], simp3511_0[0:0], simp3511_0[1:1]);
  NOR3 I391 (simp3521_0[0:0], fa3_16min_0[1:1], fa3_16min_0[2:2], fa3_16min_0[4:4]);
  INV I392 (simp3521_0[1:1], fa3_16min_0[7:7]);
  NAND2 I393 (o_0r1[16:16], simp3521_0[0:0], simp3521_0[1:1]);
  AO222 I394 (ct3__0[16:16], termt_1[16:16], termt_2[16:16], termt_1[16:16], ct3__0[15:15], termt_2[16:16], ct3__0[15:15]);
  AO222 I395 (cf3__0[16:16], termf_1[16:16], termf_2[16:16], termf_1[16:16], cf3__0[15:15], termf_2[16:16], cf3__0[15:15]);
  C3 I396 (fa3_17min_0[0:0], cf3__0[16:16], termf_2[17:17], termf_1[17:17]);
  C3 I397 (fa3_17min_0[1:1], cf3__0[16:16], termf_2[17:17], termt_1[17:17]);
  C3 I398 (fa3_17min_0[2:2], cf3__0[16:16], termt_2[17:17], termf_1[17:17]);
  C3 I399 (fa3_17min_0[3:3], cf3__0[16:16], termt_2[17:17], termt_1[17:17]);
  C3 I400 (fa3_17min_0[4:4], ct3__0[16:16], termf_2[17:17], termf_1[17:17]);
  C3 I401 (fa3_17min_0[5:5], ct3__0[16:16], termf_2[17:17], termt_1[17:17]);
  C3 I402 (fa3_17min_0[6:6], ct3__0[16:16], termt_2[17:17], termf_1[17:17]);
  C3 I403 (fa3_17min_0[7:7], ct3__0[16:16], termt_2[17:17], termt_1[17:17]);
  NOR3 I404 (simp3641_0[0:0], fa3_17min_0[0:0], fa3_17min_0[3:3], fa3_17min_0[5:5]);
  INV I405 (simp3641_0[1:1], fa3_17min_0[6:6]);
  NAND2 I406 (o_0r0[17:17], simp3641_0[0:0], simp3641_0[1:1]);
  NOR3 I407 (simp3651_0[0:0], fa3_17min_0[1:1], fa3_17min_0[2:2], fa3_17min_0[4:4]);
  INV I408 (simp3651_0[1:1], fa3_17min_0[7:7]);
  NAND2 I409 (o_0r1[17:17], simp3651_0[0:0], simp3651_0[1:1]);
  AO222 I410 (ct3__0[17:17], termt_1[17:17], termt_2[17:17], termt_1[17:17], ct3__0[16:16], termt_2[17:17], ct3__0[16:16]);
  AO222 I411 (cf3__0[17:17], termf_1[17:17], termf_2[17:17], termf_1[17:17], cf3__0[16:16], termf_2[17:17], cf3__0[16:16]);
  C3 I412 (fa3_18min_0[0:0], cf3__0[17:17], termf_2[18:18], termf_1[18:18]);
  C3 I413 (fa3_18min_0[1:1], cf3__0[17:17], termf_2[18:18], termt_1[18:18]);
  C3 I414 (fa3_18min_0[2:2], cf3__0[17:17], termt_2[18:18], termf_1[18:18]);
  C3 I415 (fa3_18min_0[3:3], cf3__0[17:17], termt_2[18:18], termt_1[18:18]);
  C3 I416 (fa3_18min_0[4:4], ct3__0[17:17], termf_2[18:18], termf_1[18:18]);
  C3 I417 (fa3_18min_0[5:5], ct3__0[17:17], termf_2[18:18], termt_1[18:18]);
  C3 I418 (fa3_18min_0[6:6], ct3__0[17:17], termt_2[18:18], termf_1[18:18]);
  C3 I419 (fa3_18min_0[7:7], ct3__0[17:17], termt_2[18:18], termt_1[18:18]);
  NOR3 I420 (simp3771_0[0:0], fa3_18min_0[0:0], fa3_18min_0[3:3], fa3_18min_0[5:5]);
  INV I421 (simp3771_0[1:1], fa3_18min_0[6:6]);
  NAND2 I422 (o_0r0[18:18], simp3771_0[0:0], simp3771_0[1:1]);
  NOR3 I423 (simp3781_0[0:0], fa3_18min_0[1:1], fa3_18min_0[2:2], fa3_18min_0[4:4]);
  INV I424 (simp3781_0[1:1], fa3_18min_0[7:7]);
  NAND2 I425 (o_0r1[18:18], simp3781_0[0:0], simp3781_0[1:1]);
  AO222 I426 (ct3__0[18:18], termt_1[18:18], termt_2[18:18], termt_1[18:18], ct3__0[17:17], termt_2[18:18], ct3__0[17:17]);
  AO222 I427 (cf3__0[18:18], termf_1[18:18], termf_2[18:18], termf_1[18:18], cf3__0[17:17], termf_2[18:18], cf3__0[17:17]);
  C3 I428 (fa3_19min_0[0:0], cf3__0[18:18], termf_2[19:19], termf_1[19:19]);
  C3 I429 (fa3_19min_0[1:1], cf3__0[18:18], termf_2[19:19], termt_1[19:19]);
  C3 I430 (fa3_19min_0[2:2], cf3__0[18:18], termt_2[19:19], termf_1[19:19]);
  C3 I431 (fa3_19min_0[3:3], cf3__0[18:18], termt_2[19:19], termt_1[19:19]);
  C3 I432 (fa3_19min_0[4:4], ct3__0[18:18], termf_2[19:19], termf_1[19:19]);
  C3 I433 (fa3_19min_0[5:5], ct3__0[18:18], termf_2[19:19], termt_1[19:19]);
  C3 I434 (fa3_19min_0[6:6], ct3__0[18:18], termt_2[19:19], termf_1[19:19]);
  C3 I435 (fa3_19min_0[7:7], ct3__0[18:18], termt_2[19:19], termt_1[19:19]);
  NOR3 I436 (simp3901_0[0:0], fa3_19min_0[0:0], fa3_19min_0[3:3], fa3_19min_0[5:5]);
  INV I437 (simp3901_0[1:1], fa3_19min_0[6:6]);
  NAND2 I438 (o_0r0[19:19], simp3901_0[0:0], simp3901_0[1:1]);
  NOR3 I439 (simp3911_0[0:0], fa3_19min_0[1:1], fa3_19min_0[2:2], fa3_19min_0[4:4]);
  INV I440 (simp3911_0[1:1], fa3_19min_0[7:7]);
  NAND2 I441 (o_0r1[19:19], simp3911_0[0:0], simp3911_0[1:1]);
  AO222 I442 (ct3__0[19:19], termt_1[19:19], termt_2[19:19], termt_1[19:19], ct3__0[18:18], termt_2[19:19], ct3__0[18:18]);
  AO222 I443 (cf3__0[19:19], termf_1[19:19], termf_2[19:19], termf_1[19:19], cf3__0[18:18], termf_2[19:19], cf3__0[18:18]);
  C3 I444 (fa3_20min_0[0:0], cf3__0[19:19], termf_2[20:20], termf_1[20:20]);
  C3 I445 (fa3_20min_0[1:1], cf3__0[19:19], termf_2[20:20], termt_1[20:20]);
  C3 I446 (fa3_20min_0[2:2], cf3__0[19:19], termt_2[20:20], termf_1[20:20]);
  C3 I447 (fa3_20min_0[3:3], cf3__0[19:19], termt_2[20:20], termt_1[20:20]);
  C3 I448 (fa3_20min_0[4:4], ct3__0[19:19], termf_2[20:20], termf_1[20:20]);
  C3 I449 (fa3_20min_0[5:5], ct3__0[19:19], termf_2[20:20], termt_1[20:20]);
  C3 I450 (fa3_20min_0[6:6], ct3__0[19:19], termt_2[20:20], termf_1[20:20]);
  C3 I451 (fa3_20min_0[7:7], ct3__0[19:19], termt_2[20:20], termt_1[20:20]);
  NOR3 I452 (simp4031_0[0:0], fa3_20min_0[0:0], fa3_20min_0[3:3], fa3_20min_0[5:5]);
  INV I453 (simp4031_0[1:1], fa3_20min_0[6:6]);
  NAND2 I454 (o_0r0[20:20], simp4031_0[0:0], simp4031_0[1:1]);
  NOR3 I455 (simp4041_0[0:0], fa3_20min_0[1:1], fa3_20min_0[2:2], fa3_20min_0[4:4]);
  INV I456 (simp4041_0[1:1], fa3_20min_0[7:7]);
  NAND2 I457 (o_0r1[20:20], simp4041_0[0:0], simp4041_0[1:1]);
  AO222 I458 (ct3__0[20:20], termt_1[20:20], termt_2[20:20], termt_1[20:20], ct3__0[19:19], termt_2[20:20], ct3__0[19:19]);
  AO222 I459 (cf3__0[20:20], termf_1[20:20], termf_2[20:20], termf_1[20:20], cf3__0[19:19], termf_2[20:20], cf3__0[19:19]);
  C3 I460 (fa3_21min_0[0:0], cf3__0[20:20], termf_2[21:21], termf_1[21:21]);
  C3 I461 (fa3_21min_0[1:1], cf3__0[20:20], termf_2[21:21], termt_1[21:21]);
  C3 I462 (fa3_21min_0[2:2], cf3__0[20:20], termt_2[21:21], termf_1[21:21]);
  C3 I463 (fa3_21min_0[3:3], cf3__0[20:20], termt_2[21:21], termt_1[21:21]);
  C3 I464 (fa3_21min_0[4:4], ct3__0[20:20], termf_2[21:21], termf_1[21:21]);
  C3 I465 (fa3_21min_0[5:5], ct3__0[20:20], termf_2[21:21], termt_1[21:21]);
  C3 I466 (fa3_21min_0[6:6], ct3__0[20:20], termt_2[21:21], termf_1[21:21]);
  C3 I467 (fa3_21min_0[7:7], ct3__0[20:20], termt_2[21:21], termt_1[21:21]);
  NOR3 I468 (simp4161_0[0:0], fa3_21min_0[0:0], fa3_21min_0[3:3], fa3_21min_0[5:5]);
  INV I469 (simp4161_0[1:1], fa3_21min_0[6:6]);
  NAND2 I470 (o_0r0[21:21], simp4161_0[0:0], simp4161_0[1:1]);
  NOR3 I471 (simp4171_0[0:0], fa3_21min_0[1:1], fa3_21min_0[2:2], fa3_21min_0[4:4]);
  INV I472 (simp4171_0[1:1], fa3_21min_0[7:7]);
  NAND2 I473 (o_0r1[21:21], simp4171_0[0:0], simp4171_0[1:1]);
  AO222 I474 (ct3__0[21:21], termt_1[21:21], termt_2[21:21], termt_1[21:21], ct3__0[20:20], termt_2[21:21], ct3__0[20:20]);
  AO222 I475 (cf3__0[21:21], termf_1[21:21], termf_2[21:21], termf_1[21:21], cf3__0[20:20], termf_2[21:21], cf3__0[20:20]);
  C3 I476 (fa3_22min_0[0:0], cf3__0[21:21], termf_2[22:22], termf_1[22:22]);
  C3 I477 (fa3_22min_0[1:1], cf3__0[21:21], termf_2[22:22], termt_1[22:22]);
  C3 I478 (fa3_22min_0[2:2], cf3__0[21:21], termt_2[22:22], termf_1[22:22]);
  C3 I479 (fa3_22min_0[3:3], cf3__0[21:21], termt_2[22:22], termt_1[22:22]);
  C3 I480 (fa3_22min_0[4:4], ct3__0[21:21], termf_2[22:22], termf_1[22:22]);
  C3 I481 (fa3_22min_0[5:5], ct3__0[21:21], termf_2[22:22], termt_1[22:22]);
  C3 I482 (fa3_22min_0[6:6], ct3__0[21:21], termt_2[22:22], termf_1[22:22]);
  C3 I483 (fa3_22min_0[7:7], ct3__0[21:21], termt_2[22:22], termt_1[22:22]);
  NOR3 I484 (simp4291_0[0:0], fa3_22min_0[0:0], fa3_22min_0[3:3], fa3_22min_0[5:5]);
  INV I485 (simp4291_0[1:1], fa3_22min_0[6:6]);
  NAND2 I486 (o_0r0[22:22], simp4291_0[0:0], simp4291_0[1:1]);
  NOR3 I487 (simp4301_0[0:0], fa3_22min_0[1:1], fa3_22min_0[2:2], fa3_22min_0[4:4]);
  INV I488 (simp4301_0[1:1], fa3_22min_0[7:7]);
  NAND2 I489 (o_0r1[22:22], simp4301_0[0:0], simp4301_0[1:1]);
  AO222 I490 (ct3__0[22:22], termt_1[22:22], termt_2[22:22], termt_1[22:22], ct3__0[21:21], termt_2[22:22], ct3__0[21:21]);
  AO222 I491 (cf3__0[22:22], termf_1[22:22], termf_2[22:22], termf_1[22:22], cf3__0[21:21], termf_2[22:22], cf3__0[21:21]);
  C3 I492 (fa3_23min_0[0:0], cf3__0[22:22], termf_2[23:23], termf_1[23:23]);
  C3 I493 (fa3_23min_0[1:1], cf3__0[22:22], termf_2[23:23], termt_1[23:23]);
  C3 I494 (fa3_23min_0[2:2], cf3__0[22:22], termt_2[23:23], termf_1[23:23]);
  C3 I495 (fa3_23min_0[3:3], cf3__0[22:22], termt_2[23:23], termt_1[23:23]);
  C3 I496 (fa3_23min_0[4:4], ct3__0[22:22], termf_2[23:23], termf_1[23:23]);
  C3 I497 (fa3_23min_0[5:5], ct3__0[22:22], termf_2[23:23], termt_1[23:23]);
  C3 I498 (fa3_23min_0[6:6], ct3__0[22:22], termt_2[23:23], termf_1[23:23]);
  C3 I499 (fa3_23min_0[7:7], ct3__0[22:22], termt_2[23:23], termt_1[23:23]);
  NOR3 I500 (simp4421_0[0:0], fa3_23min_0[0:0], fa3_23min_0[3:3], fa3_23min_0[5:5]);
  INV I501 (simp4421_0[1:1], fa3_23min_0[6:6]);
  NAND2 I502 (o_0r0[23:23], simp4421_0[0:0], simp4421_0[1:1]);
  NOR3 I503 (simp4431_0[0:0], fa3_23min_0[1:1], fa3_23min_0[2:2], fa3_23min_0[4:4]);
  INV I504 (simp4431_0[1:1], fa3_23min_0[7:7]);
  NAND2 I505 (o_0r1[23:23], simp4431_0[0:0], simp4431_0[1:1]);
  AO222 I506 (ct3__0[23:23], termt_1[23:23], termt_2[23:23], termt_1[23:23], ct3__0[22:22], termt_2[23:23], ct3__0[22:22]);
  AO222 I507 (cf3__0[23:23], termf_1[23:23], termf_2[23:23], termf_1[23:23], cf3__0[22:22], termf_2[23:23], cf3__0[22:22]);
  C3 I508 (fa3_24min_0[0:0], cf3__0[23:23], termf_2[24:24], termf_1[24:24]);
  C3 I509 (fa3_24min_0[1:1], cf3__0[23:23], termf_2[24:24], termt_1[24:24]);
  C3 I510 (fa3_24min_0[2:2], cf3__0[23:23], termt_2[24:24], termf_1[24:24]);
  C3 I511 (fa3_24min_0[3:3], cf3__0[23:23], termt_2[24:24], termt_1[24:24]);
  C3 I512 (fa3_24min_0[4:4], ct3__0[23:23], termf_2[24:24], termf_1[24:24]);
  C3 I513 (fa3_24min_0[5:5], ct3__0[23:23], termf_2[24:24], termt_1[24:24]);
  C3 I514 (fa3_24min_0[6:6], ct3__0[23:23], termt_2[24:24], termf_1[24:24]);
  C3 I515 (fa3_24min_0[7:7], ct3__0[23:23], termt_2[24:24], termt_1[24:24]);
  NOR3 I516 (simp4551_0[0:0], fa3_24min_0[0:0], fa3_24min_0[3:3], fa3_24min_0[5:5]);
  INV I517 (simp4551_0[1:1], fa3_24min_0[6:6]);
  NAND2 I518 (o_0r0[24:24], simp4551_0[0:0], simp4551_0[1:1]);
  NOR3 I519 (simp4561_0[0:0], fa3_24min_0[1:1], fa3_24min_0[2:2], fa3_24min_0[4:4]);
  INV I520 (simp4561_0[1:1], fa3_24min_0[7:7]);
  NAND2 I521 (o_0r1[24:24], simp4561_0[0:0], simp4561_0[1:1]);
  AO222 I522 (ct3__0[24:24], termt_1[24:24], termt_2[24:24], termt_1[24:24], ct3__0[23:23], termt_2[24:24], ct3__0[23:23]);
  AO222 I523 (cf3__0[24:24], termf_1[24:24], termf_2[24:24], termf_1[24:24], cf3__0[23:23], termf_2[24:24], cf3__0[23:23]);
  C3 I524 (fa3_25min_0[0:0], cf3__0[24:24], termf_2[25:25], termf_1[25:25]);
  C3 I525 (fa3_25min_0[1:1], cf3__0[24:24], termf_2[25:25], termt_1[25:25]);
  C3 I526 (fa3_25min_0[2:2], cf3__0[24:24], termt_2[25:25], termf_1[25:25]);
  C3 I527 (fa3_25min_0[3:3], cf3__0[24:24], termt_2[25:25], termt_1[25:25]);
  C3 I528 (fa3_25min_0[4:4], ct3__0[24:24], termf_2[25:25], termf_1[25:25]);
  C3 I529 (fa3_25min_0[5:5], ct3__0[24:24], termf_2[25:25], termt_1[25:25]);
  C3 I530 (fa3_25min_0[6:6], ct3__0[24:24], termt_2[25:25], termf_1[25:25]);
  C3 I531 (fa3_25min_0[7:7], ct3__0[24:24], termt_2[25:25], termt_1[25:25]);
  NOR3 I532 (simp4681_0[0:0], fa3_25min_0[0:0], fa3_25min_0[3:3], fa3_25min_0[5:5]);
  INV I533 (simp4681_0[1:1], fa3_25min_0[6:6]);
  NAND2 I534 (o_0r0[25:25], simp4681_0[0:0], simp4681_0[1:1]);
  NOR3 I535 (simp4691_0[0:0], fa3_25min_0[1:1], fa3_25min_0[2:2], fa3_25min_0[4:4]);
  INV I536 (simp4691_0[1:1], fa3_25min_0[7:7]);
  NAND2 I537 (o_0r1[25:25], simp4691_0[0:0], simp4691_0[1:1]);
  AO222 I538 (ct3__0[25:25], termt_1[25:25], termt_2[25:25], termt_1[25:25], ct3__0[24:24], termt_2[25:25], ct3__0[24:24]);
  AO222 I539 (cf3__0[25:25], termf_1[25:25], termf_2[25:25], termf_1[25:25], cf3__0[24:24], termf_2[25:25], cf3__0[24:24]);
  C3 I540 (fa3_26min_0[0:0], cf3__0[25:25], termf_2[26:26], termf_1[26:26]);
  C3 I541 (fa3_26min_0[1:1], cf3__0[25:25], termf_2[26:26], termt_1[26:26]);
  C3 I542 (fa3_26min_0[2:2], cf3__0[25:25], termt_2[26:26], termf_1[26:26]);
  C3 I543 (fa3_26min_0[3:3], cf3__0[25:25], termt_2[26:26], termt_1[26:26]);
  C3 I544 (fa3_26min_0[4:4], ct3__0[25:25], termf_2[26:26], termf_1[26:26]);
  C3 I545 (fa3_26min_0[5:5], ct3__0[25:25], termf_2[26:26], termt_1[26:26]);
  C3 I546 (fa3_26min_0[6:6], ct3__0[25:25], termt_2[26:26], termf_1[26:26]);
  C3 I547 (fa3_26min_0[7:7], ct3__0[25:25], termt_2[26:26], termt_1[26:26]);
  NOR3 I548 (simp4811_0[0:0], fa3_26min_0[0:0], fa3_26min_0[3:3], fa3_26min_0[5:5]);
  INV I549 (simp4811_0[1:1], fa3_26min_0[6:6]);
  NAND2 I550 (o_0r0[26:26], simp4811_0[0:0], simp4811_0[1:1]);
  NOR3 I551 (simp4821_0[0:0], fa3_26min_0[1:1], fa3_26min_0[2:2], fa3_26min_0[4:4]);
  INV I552 (simp4821_0[1:1], fa3_26min_0[7:7]);
  NAND2 I553 (o_0r1[26:26], simp4821_0[0:0], simp4821_0[1:1]);
  AO222 I554 (ct3__0[26:26], termt_1[26:26], termt_2[26:26], termt_1[26:26], ct3__0[25:25], termt_2[26:26], ct3__0[25:25]);
  AO222 I555 (cf3__0[26:26], termf_1[26:26], termf_2[26:26], termf_1[26:26], cf3__0[25:25], termf_2[26:26], cf3__0[25:25]);
  C3 I556 (fa3_27min_0[0:0], cf3__0[26:26], termf_2[27:27], termf_1[27:27]);
  C3 I557 (fa3_27min_0[1:1], cf3__0[26:26], termf_2[27:27], termt_1[27:27]);
  C3 I558 (fa3_27min_0[2:2], cf3__0[26:26], termt_2[27:27], termf_1[27:27]);
  C3 I559 (fa3_27min_0[3:3], cf3__0[26:26], termt_2[27:27], termt_1[27:27]);
  C3 I560 (fa3_27min_0[4:4], ct3__0[26:26], termf_2[27:27], termf_1[27:27]);
  C3 I561 (fa3_27min_0[5:5], ct3__0[26:26], termf_2[27:27], termt_1[27:27]);
  C3 I562 (fa3_27min_0[6:6], ct3__0[26:26], termt_2[27:27], termf_1[27:27]);
  C3 I563 (fa3_27min_0[7:7], ct3__0[26:26], termt_2[27:27], termt_1[27:27]);
  NOR3 I564 (simp4941_0[0:0], fa3_27min_0[0:0], fa3_27min_0[3:3], fa3_27min_0[5:5]);
  INV I565 (simp4941_0[1:1], fa3_27min_0[6:6]);
  NAND2 I566 (o_0r0[27:27], simp4941_0[0:0], simp4941_0[1:1]);
  NOR3 I567 (simp4951_0[0:0], fa3_27min_0[1:1], fa3_27min_0[2:2], fa3_27min_0[4:4]);
  INV I568 (simp4951_0[1:1], fa3_27min_0[7:7]);
  NAND2 I569 (o_0r1[27:27], simp4951_0[0:0], simp4951_0[1:1]);
  AO222 I570 (ct3__0[27:27], termt_1[27:27], termt_2[27:27], termt_1[27:27], ct3__0[26:26], termt_2[27:27], ct3__0[26:26]);
  AO222 I571 (cf3__0[27:27], termf_1[27:27], termf_2[27:27], termf_1[27:27], cf3__0[26:26], termf_2[27:27], cf3__0[26:26]);
  C3 I572 (fa3_28min_0[0:0], cf3__0[27:27], termf_2[28:28], termf_1[28:28]);
  C3 I573 (fa3_28min_0[1:1], cf3__0[27:27], termf_2[28:28], termt_1[28:28]);
  C3 I574 (fa3_28min_0[2:2], cf3__0[27:27], termt_2[28:28], termf_1[28:28]);
  C3 I575 (fa3_28min_0[3:3], cf3__0[27:27], termt_2[28:28], termt_1[28:28]);
  C3 I576 (fa3_28min_0[4:4], ct3__0[27:27], termf_2[28:28], termf_1[28:28]);
  C3 I577 (fa3_28min_0[5:5], ct3__0[27:27], termf_2[28:28], termt_1[28:28]);
  C3 I578 (fa3_28min_0[6:6], ct3__0[27:27], termt_2[28:28], termf_1[28:28]);
  C3 I579 (fa3_28min_0[7:7], ct3__0[27:27], termt_2[28:28], termt_1[28:28]);
  NOR3 I580 (simp5071_0[0:0], fa3_28min_0[0:0], fa3_28min_0[3:3], fa3_28min_0[5:5]);
  INV I581 (simp5071_0[1:1], fa3_28min_0[6:6]);
  NAND2 I582 (o_0r0[28:28], simp5071_0[0:0], simp5071_0[1:1]);
  NOR3 I583 (simp5081_0[0:0], fa3_28min_0[1:1], fa3_28min_0[2:2], fa3_28min_0[4:4]);
  INV I584 (simp5081_0[1:1], fa3_28min_0[7:7]);
  NAND2 I585 (o_0r1[28:28], simp5081_0[0:0], simp5081_0[1:1]);
  AO222 I586 (ct3__0[28:28], termt_1[28:28], termt_2[28:28], termt_1[28:28], ct3__0[27:27], termt_2[28:28], ct3__0[27:27]);
  AO222 I587 (cf3__0[28:28], termf_1[28:28], termf_2[28:28], termf_1[28:28], cf3__0[27:27], termf_2[28:28], cf3__0[27:27]);
  C3 I588 (fa3_29min_0[0:0], cf3__0[28:28], termf_2[29:29], termf_1[29:29]);
  C3 I589 (fa3_29min_0[1:1], cf3__0[28:28], termf_2[29:29], termt_1[29:29]);
  C3 I590 (fa3_29min_0[2:2], cf3__0[28:28], termt_2[29:29], termf_1[29:29]);
  C3 I591 (fa3_29min_0[3:3], cf3__0[28:28], termt_2[29:29], termt_1[29:29]);
  C3 I592 (fa3_29min_0[4:4], ct3__0[28:28], termf_2[29:29], termf_1[29:29]);
  C3 I593 (fa3_29min_0[5:5], ct3__0[28:28], termf_2[29:29], termt_1[29:29]);
  C3 I594 (fa3_29min_0[6:6], ct3__0[28:28], termt_2[29:29], termf_1[29:29]);
  C3 I595 (fa3_29min_0[7:7], ct3__0[28:28], termt_2[29:29], termt_1[29:29]);
  NOR3 I596 (simp5201_0[0:0], fa3_29min_0[0:0], fa3_29min_0[3:3], fa3_29min_0[5:5]);
  INV I597 (simp5201_0[1:1], fa3_29min_0[6:6]);
  NAND2 I598 (o_0r0[29:29], simp5201_0[0:0], simp5201_0[1:1]);
  NOR3 I599 (simp5211_0[0:0], fa3_29min_0[1:1], fa3_29min_0[2:2], fa3_29min_0[4:4]);
  INV I600 (simp5211_0[1:1], fa3_29min_0[7:7]);
  NAND2 I601 (o_0r1[29:29], simp5211_0[0:0], simp5211_0[1:1]);
  AO222 I602 (ct3__0[29:29], termt_1[29:29], termt_2[29:29], termt_1[29:29], ct3__0[28:28], termt_2[29:29], ct3__0[28:28]);
  AO222 I603 (cf3__0[29:29], termf_1[29:29], termf_2[29:29], termf_1[29:29], cf3__0[28:28], termf_2[29:29], cf3__0[28:28]);
  C3 I604 (fa3_30min_0[0:0], cf3__0[29:29], termf_2[30:30], termf_1[30:30]);
  C3 I605 (fa3_30min_0[1:1], cf3__0[29:29], termf_2[30:30], termt_1[30:30]);
  C3 I606 (fa3_30min_0[2:2], cf3__0[29:29], termt_2[30:30], termf_1[30:30]);
  C3 I607 (fa3_30min_0[3:3], cf3__0[29:29], termt_2[30:30], termt_1[30:30]);
  C3 I608 (fa3_30min_0[4:4], ct3__0[29:29], termf_2[30:30], termf_1[30:30]);
  C3 I609 (fa3_30min_0[5:5], ct3__0[29:29], termf_2[30:30], termt_1[30:30]);
  C3 I610 (fa3_30min_0[6:6], ct3__0[29:29], termt_2[30:30], termf_1[30:30]);
  C3 I611 (fa3_30min_0[7:7], ct3__0[29:29], termt_2[30:30], termt_1[30:30]);
  NOR3 I612 (simp5331_0[0:0], fa3_30min_0[0:0], fa3_30min_0[3:3], fa3_30min_0[5:5]);
  INV I613 (simp5331_0[1:1], fa3_30min_0[6:6]);
  NAND2 I614 (o_0r0[30:30], simp5331_0[0:0], simp5331_0[1:1]);
  NOR3 I615 (simp5341_0[0:0], fa3_30min_0[1:1], fa3_30min_0[2:2], fa3_30min_0[4:4]);
  INV I616 (simp5341_0[1:1], fa3_30min_0[7:7]);
  NAND2 I617 (o_0r1[30:30], simp5341_0[0:0], simp5341_0[1:1]);
  AO222 I618 (ct3__0[30:30], termt_1[30:30], termt_2[30:30], termt_1[30:30], ct3__0[29:29], termt_2[30:30], ct3__0[29:29]);
  AO222 I619 (cf3__0[30:30], termf_1[30:30], termf_2[30:30], termf_1[30:30], cf3__0[29:29], termf_2[30:30], cf3__0[29:29]);
  C3 I620 (fa3_31min_0[0:0], cf3__0[30:30], termf_2[31:31], termf_1[31:31]);
  C3 I621 (fa3_31min_0[1:1], cf3__0[30:30], termf_2[31:31], termt_1[31:31]);
  C3 I622 (fa3_31min_0[2:2], cf3__0[30:30], termt_2[31:31], termf_1[31:31]);
  C3 I623 (fa3_31min_0[3:3], cf3__0[30:30], termt_2[31:31], termt_1[31:31]);
  C3 I624 (fa3_31min_0[4:4], ct3__0[30:30], termf_2[31:31], termf_1[31:31]);
  C3 I625 (fa3_31min_0[5:5], ct3__0[30:30], termf_2[31:31], termt_1[31:31]);
  C3 I626 (fa3_31min_0[6:6], ct3__0[30:30], termt_2[31:31], termf_1[31:31]);
  C3 I627 (fa3_31min_0[7:7], ct3__0[30:30], termt_2[31:31], termt_1[31:31]);
  NOR3 I628 (simp5461_0[0:0], fa3_31min_0[0:0], fa3_31min_0[3:3], fa3_31min_0[5:5]);
  INV I629 (simp5461_0[1:1], fa3_31min_0[6:6]);
  NAND2 I630 (o_0r0[31:31], simp5461_0[0:0], simp5461_0[1:1]);
  NOR3 I631 (simp5471_0[0:0], fa3_31min_0[1:1], fa3_31min_0[2:2], fa3_31min_0[4:4]);
  INV I632 (simp5471_0[1:1], fa3_31min_0[7:7]);
  NAND2 I633 (o_0r1[31:31], simp5471_0[0:0], simp5471_0[1:1]);
  AO222 I634 (ct3__0[31:31], termt_1[31:31], termt_2[31:31], termt_1[31:31], ct3__0[30:30], termt_2[31:31], ct3__0[30:30]);
  AO222 I635 (cf3__0[31:31], termf_1[31:31], termf_2[31:31], termf_1[31:31], cf3__0[30:30], termf_2[31:31], cf3__0[30:30]);
  C3 I636 (fa3_32min_0[0:0], cf3__0[31:31], termf_2[32:32], termf_1[32:32]);
  C3 I637 (fa3_32min_0[1:1], cf3__0[31:31], termf_2[32:32], termt_1[32:32]);
  C3 I638 (fa3_32min_0[2:2], cf3__0[31:31], termt_2[32:32], termf_1[32:32]);
  C3 I639 (fa3_32min_0[3:3], cf3__0[31:31], termt_2[32:32], termt_1[32:32]);
  C3 I640 (fa3_32min_0[4:4], ct3__0[31:31], termf_2[32:32], termf_1[32:32]);
  C3 I641 (fa3_32min_0[5:5], ct3__0[31:31], termf_2[32:32], termt_1[32:32]);
  C3 I642 (fa3_32min_0[6:6], ct3__0[31:31], termt_2[32:32], termf_1[32:32]);
  C3 I643 (fa3_32min_0[7:7], ct3__0[31:31], termt_2[32:32], termt_1[32:32]);
  NOR3 I644 (simp5591_0[0:0], fa3_32min_0[0:0], fa3_32min_0[3:3], fa3_32min_0[5:5]);
  INV I645 (simp5591_0[1:1], fa3_32min_0[6:6]);
  NAND2 I646 (o_0r0[32:32], simp5591_0[0:0], simp5591_0[1:1]);
  NOR3 I647 (simp5601_0[0:0], fa3_32min_0[1:1], fa3_32min_0[2:2], fa3_32min_0[4:4]);
  INV I648 (simp5601_0[1:1], fa3_32min_0[7:7]);
  NAND2 I649 (o_0r1[32:32], simp5601_0[0:0], simp5601_0[1:1]);
  AO222 I650 (ct3__0[32:32], termt_1[32:32], termt_2[32:32], termt_1[32:32], ct3__0[31:31], termt_2[32:32], ct3__0[31:31]);
  AO222 I651 (cf3__0[32:32], termf_1[32:32], termf_2[32:32], termf_1[32:32], cf3__0[31:31], termf_2[32:32], cf3__0[31:31]);
  BUFF I652 (i_0a, o_0a);
endmodule

// tkf33mo0w0_o0w32 TeakF [0,0] [One 33,Many [0,32]]
module tkf33mo0w0_o0w32 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire comp_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0, i_0r0[32:32], i_0r1[32:32]);
  BUFF I2 (ucomplete_0, comp_0);
  C2 I3 (acomplete_0, ucomplete_0, icomplete_0);
  C2 I4 (o_1r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I5 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I6 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I7 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I8 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I9 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I10 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I11 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I12 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I13 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I14 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I15 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I16 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I17 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I18 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I19 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I20 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I21 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I22 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I23 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I24 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I25 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I26 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I27 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I28 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I29 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I30 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I31 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I32 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I33 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I34 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I35 (o_1r0[31:31], i_0r0[31:31]);
  C2 I36 (o_1r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I37 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I38 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I39 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I40 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I41 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I42 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I43 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I44 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I45 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I46 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I47 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I48 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I49 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I50 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I51 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I52 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I53 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I54 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I55 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I56 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I57 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I58 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I59 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I60 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I61 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I62 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I63 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I64 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I65 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I66 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I67 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I68 (o_0r, icomplete_0);
  C3 I69 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkf0mo0w0_o0w0 TeakF [0,0] [One 0,Many [0,0]]
module tkf0mo0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  C2 I2 (i_0a, o_0a, o_1a);
endmodule

// tkm3x0b TeakM [Many [0,0,0],One 0]
module tkm3x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  NOR2 I3 (nchosen_0, o_0r, o_0a);
  OR3 I4 (o_0r, choice_0, choice_1, choice_2);
  C2R I5 (i_0a, choice_0, o_0a, reset);
  C2R I6 (i_1a, choice_1, o_0a, reset);
  C2R I7 (i_2a, choice_2, o_0a, reset);
endmodule

// tkm3x3b TeakM [Many [3,3,3],One 3]
module tkm3x3b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  input [2:0] i_2r0;
  input [2:0] i_2r1;
  output i_2a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire [2:0] gfint_0;
  wire [2:0] gfint_1;
  wire [2:0] gfint_2;
  wire [2:0] gtint_0;
  wire [2:0] gtint_1;
  wire [2:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [2:0] comp0_0;
  wire [2:0] comp1_0;
  wire [2:0] comp2_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  OR3 I3 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I4 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  OR3 I5 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  AND2 I6 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I7 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I8 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I9 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I10 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I11 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I12 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I13 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I14 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I15 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I16 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I17 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I18 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I19 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I20 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I21 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I22 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I23 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  OR2 I24 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I27 (icomp_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  OR2 I28 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I29 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I30 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  C3 I31 (icomp_1, comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  OR2 I32 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I33 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I34 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  C3 I35 (icomp_2, comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C2R I36 (choice_0, icomp_0, nchosen_0, reset);
  C2R I37 (choice_1, icomp_1, nchosen_0, reset);
  C2R I38 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I39 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I40 (nchosen_0, anychoice_0, o_0a);
  C2R I41 (i_0a, choice_0, o_0a, reset);
  C2R I42 (i_1a, choice_1, o_0a, reset);
  C2R I43 (i_2a, choice_2, o_0a, reset);
endmodule

// tko0m3_1nm3b1 TeakO [
//     (1,TeakOConstant 3 1)] [One 0,One 3]
module tko0m3_1nm3b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  GND I4 (o_0r1[1:1]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b2 TeakO [
//     (1,TeakOConstant 3 2)] [One 0,One 3]
module tko0m3_1nm3b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  GND I4 (o_0r1[0:0]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b4 TeakO [
//     (1,TeakOConstant 3 4)] [One 0,One 3]
module tko0m3_1nm3b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  GND I4 (o_0r1[0:0]);
  GND I5 (o_0r1[1:1]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tkj3m0_3 TeakJ [Many [0,3],One 3]
module tkj3m0_3 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joint_0[0:0], i_1r1[0:0]);
  BUFF I4 (joint_0[1:1], i_1r1[1:1]);
  BUFF I5 (joint_0[2:2], i_1r1[2:2]);
  BUFF I6 (icomplete_0, i_0r);
  C2 I7 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I8 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I9 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I10 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I11 (o_0r1[1:1], joint_0[1:1]);
  BUFF I12 (o_0r1[2:2], joint_0[2:2]);
  BUFF I13 (i_0a, o_0a);
  BUFF I14 (i_1a, o_0a);
endmodule

// tks3_o0w3_1o0w0_2o0w0_4o0w0 TeakS (0+:3) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0)] [One 3,Many [0,
//   0,0]]
module tks3_o0w3_1o0w0_2o0w0_4o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [2:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I11 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I12 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I13 (o_0r, gsel_0);
  BUFF I14 (o_1r, gsel_1);
  BUFF I15 (o_2r, gsel_2);
  OR3 I16 (oack_0, o_0a, o_1a, o_2a);
  C2 I17 (i_0a, oack_0, icomplete_0);
endmodule

// tkvneg3_wo0w3_ro0w3o0w3o0w3 TeakV "neg" 3 [] [0] [0,0,0] [Many [3],Many [0],Many [0,0,0],Many [3,3,3
//   ]]
module tkvneg3_wo0w3_ro0w3o0w3o0w3 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [2:0] wg_0r0;
  input [2:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [2:0] rd_0r0;
  output [2:0] rd_0r1;
  input rd_0a;
  output [2:0] rd_1r0;
  output [2:0] rd_1r1;
  input rd_1a;
  output [2:0] rd_2r0;
  output [2:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [2:0] wf_0;
  wire [2:0] wt_0;
  wire [2:0] df_0;
  wire [2:0] dt_0;
  wire wc_0;
  wire [2:0] wacks_0;
  wire [2:0] wenr_0;
  wire [2:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [2:0] drlgf_0;
  wire [2:0] drlgt_0;
  wire [2:0] comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [2:0] conwgit_0;
  wire [2:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp591_0;
  wire [1:0] simp781_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I5 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I6 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I7 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I8 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I9 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  NOR2 I10 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I11 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I12 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR3 I13 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I14 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I15 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  AO22 I16 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I17 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I18 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  OR2 I19 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I20 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I21 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  C3 I22 (wc_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  AND2 I23 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I24 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I25 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I26 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I27 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I28 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  BUFF I29 (conwigc_0, wc_0);
  AO22 I30 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I31 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I32 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I33 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I34 (wenr_0[0:0], wc_0);
  BUFF I35 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I36 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I37 (wenr_0[1:1], wc_0);
  BUFF I38 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I39 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I40 (wenr_0[2:2], wc_0);
  C3 I41 (simp591_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  BUFF I42 (simp591_0[1:1], wacks_0[2:2]);
  C2 I43 (wd_0r, simp591_0[0:0], simp591_0[1:1]);
  AND2 I44 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I45 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I46 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I47 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I48 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I49 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I50 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I51 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I52 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I53 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I54 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I55 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I56 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I57 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I58 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I59 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I60 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I61 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  NOR3 I62 (simp781_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I63 (simp781_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I64 (anyread_0, simp781_0[0:0], simp781_0[1:1]);
  BUFF I65 (wg_0a, wd_0a);
  BUFF I66 (rg_0a, rd_0a);
  BUFF I67 (rg_1a, rd_1a);
  BUFF I68 (rg_2a, rd_2a);
endmodule

// tkm3x32b TeakM [Many [32,32,32],One 32]
module tkm3x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [31:0] comp0_0;
  wire [10:0] simp3031_0;
  wire [3:0] simp3032_0;
  wire [1:0] simp3033_0;
  wire [31:0] comp1_0;
  wire [10:0] simp3371_0;
  wire [3:0] simp3372_0;
  wire [1:0] simp3373_0;
  wire [31:0] comp2_0;
  wire [10:0] simp3711_0;
  wire [3:0] simp3712_0;
  wire [1:0] simp3713_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  OR3 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  OR3 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  OR3 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  OR3 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  OR3 I7 (o_0r0[7:7], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  OR3 I8 (o_0r0[8:8], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  OR3 I9 (o_0r0[9:9], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  OR3 I10 (o_0r0[10:10], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  OR3 I11 (o_0r0[11:11], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  OR3 I12 (o_0r0[12:12], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  OR3 I13 (o_0r0[13:13], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  OR3 I14 (o_0r0[14:14], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  OR3 I15 (o_0r0[15:15], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  OR3 I16 (o_0r0[16:16], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  OR3 I17 (o_0r0[17:17], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  OR3 I18 (o_0r0[18:18], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  OR3 I19 (o_0r0[19:19], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  OR3 I20 (o_0r0[20:20], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  OR3 I21 (o_0r0[21:21], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  OR3 I22 (o_0r0[22:22], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  OR3 I23 (o_0r0[23:23], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  OR3 I24 (o_0r0[24:24], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  OR3 I25 (o_0r0[25:25], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  OR3 I26 (o_0r0[26:26], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  OR3 I27 (o_0r0[27:27], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  OR3 I28 (o_0r0[28:28], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  OR3 I29 (o_0r0[29:29], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  OR3 I30 (o_0r0[30:30], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  OR3 I31 (o_0r0[31:31], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  OR3 I32 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I33 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  OR3 I34 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  OR3 I35 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  OR3 I36 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  OR3 I37 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  OR3 I38 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  OR3 I39 (o_0r1[7:7], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  OR3 I40 (o_0r1[8:8], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  OR3 I41 (o_0r1[9:9], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  OR3 I42 (o_0r1[10:10], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  OR3 I43 (o_0r1[11:11], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  OR3 I44 (o_0r1[12:12], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  OR3 I45 (o_0r1[13:13], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  OR3 I46 (o_0r1[14:14], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  OR3 I47 (o_0r1[15:15], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  OR3 I48 (o_0r1[16:16], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  OR3 I49 (o_0r1[17:17], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  OR3 I50 (o_0r1[18:18], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  OR3 I51 (o_0r1[19:19], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  OR3 I52 (o_0r1[20:20], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  OR3 I53 (o_0r1[21:21], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  OR3 I54 (o_0r1[22:22], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  OR3 I55 (o_0r1[23:23], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  OR3 I56 (o_0r1[24:24], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  OR3 I57 (o_0r1[25:25], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  OR3 I58 (o_0r1[26:26], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  OR3 I59 (o_0r1[27:27], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  OR3 I60 (o_0r1[28:28], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  OR3 I61 (o_0r1[29:29], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  OR3 I62 (o_0r1[30:30], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  OR3 I63 (o_0r1[31:31], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  AND2 I64 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I65 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I66 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I67 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I68 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I69 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I70 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I71 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I72 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I73 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I74 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I75 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I76 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I77 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I78 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I79 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I80 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I81 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I82 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I83 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I84 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I85 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I86 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I87 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I88 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I89 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I90 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I91 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I92 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I93 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I94 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I95 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I96 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I97 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I98 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I99 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I100 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I101 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I102 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I103 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I104 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I105 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I106 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I107 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I108 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I109 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I110 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I111 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I112 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I113 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I114 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I115 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I116 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I117 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I118 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I119 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I120 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I121 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I122 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I123 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I124 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I125 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I126 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I127 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I128 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I129 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I130 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I131 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I132 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I133 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I134 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I135 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I136 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I137 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I138 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I139 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I140 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I141 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I142 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I143 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I144 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I145 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I146 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I147 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I148 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I149 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I150 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I151 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I152 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I153 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I154 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I155 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I156 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I157 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I158 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I159 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I160 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I161 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I162 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I163 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I164 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I165 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I166 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I167 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I168 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I169 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I170 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I171 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I172 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I173 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I174 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I175 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I176 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I177 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I178 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I179 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I180 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I181 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I182 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I183 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I184 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I185 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I186 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I187 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I188 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I189 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I190 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I191 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I192 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I193 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I194 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I195 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I196 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I197 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I198 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I199 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I200 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I201 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I202 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I203 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I204 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I205 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I206 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I207 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I208 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I209 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I210 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I211 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I212 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I213 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I214 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I215 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I216 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I217 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I218 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I219 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I220 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I221 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I222 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I223 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I224 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I225 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I226 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I227 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I228 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I229 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I230 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I231 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I232 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I233 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I234 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I235 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I236 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I237 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I238 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I239 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I240 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I241 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I242 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I243 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I244 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I245 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I246 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I247 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I248 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I249 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I250 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I251 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I252 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I253 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I254 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I255 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  OR2 I256 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I257 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I258 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I259 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I260 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I261 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I262 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I263 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I264 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I265 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I266 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I267 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I268 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I269 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I270 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I271 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I272 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I273 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I274 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I275 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I276 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I277 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I278 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I279 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I280 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I281 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I282 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I283 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I284 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I285 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I286 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I287 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I288 (simp3031_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I289 (simp3031_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I290 (simp3031_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I291 (simp3031_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I292 (simp3031_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I293 (simp3031_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I294 (simp3031_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I295 (simp3031_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I296 (simp3031_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I297 (simp3031_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I298 (simp3031_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I299 (simp3032_0[0:0], simp3031_0[0:0], simp3031_0[1:1], simp3031_0[2:2]);
  C3 I300 (simp3032_0[1:1], simp3031_0[3:3], simp3031_0[4:4], simp3031_0[5:5]);
  C3 I301 (simp3032_0[2:2], simp3031_0[6:6], simp3031_0[7:7], simp3031_0[8:8]);
  C2 I302 (simp3032_0[3:3], simp3031_0[9:9], simp3031_0[10:10]);
  C3 I303 (simp3033_0[0:0], simp3032_0[0:0], simp3032_0[1:1], simp3032_0[2:2]);
  BUFF I304 (simp3033_0[1:1], simp3032_0[3:3]);
  C2 I305 (icomp_0, simp3033_0[0:0], simp3033_0[1:1]);
  OR2 I306 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I307 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I308 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I309 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I310 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I311 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I312 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I313 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I314 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I315 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I316 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I317 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I318 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I319 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I320 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I321 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I322 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I323 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I324 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I325 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I326 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I327 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I328 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I329 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I330 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I331 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I332 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I333 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I334 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I335 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I336 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I337 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I338 (simp3371_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I339 (simp3371_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I340 (simp3371_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I341 (simp3371_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I342 (simp3371_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I343 (simp3371_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I344 (simp3371_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I345 (simp3371_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I346 (simp3371_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I347 (simp3371_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I348 (simp3371_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I349 (simp3372_0[0:0], simp3371_0[0:0], simp3371_0[1:1], simp3371_0[2:2]);
  C3 I350 (simp3372_0[1:1], simp3371_0[3:3], simp3371_0[4:4], simp3371_0[5:5]);
  C3 I351 (simp3372_0[2:2], simp3371_0[6:6], simp3371_0[7:7], simp3371_0[8:8]);
  C2 I352 (simp3372_0[3:3], simp3371_0[9:9], simp3371_0[10:10]);
  C3 I353 (simp3373_0[0:0], simp3372_0[0:0], simp3372_0[1:1], simp3372_0[2:2]);
  BUFF I354 (simp3373_0[1:1], simp3372_0[3:3]);
  C2 I355 (icomp_1, simp3373_0[0:0], simp3373_0[1:1]);
  OR2 I356 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I357 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I358 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I359 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I360 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I361 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I362 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I363 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I364 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I365 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I366 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I367 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I368 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I369 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I370 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I371 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I372 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I373 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I374 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I375 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I376 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I377 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I378 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I379 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I380 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I381 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I382 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I383 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I384 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I385 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I386 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I387 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  C3 I388 (simp3711_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I389 (simp3711_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I390 (simp3711_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I391 (simp3711_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I392 (simp3711_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I393 (simp3711_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I394 (simp3711_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I395 (simp3711_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I396 (simp3711_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I397 (simp3711_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C2 I398 (simp3711_0[10:10], comp2_0[30:30], comp2_0[31:31]);
  C3 I399 (simp3712_0[0:0], simp3711_0[0:0], simp3711_0[1:1], simp3711_0[2:2]);
  C3 I400 (simp3712_0[1:1], simp3711_0[3:3], simp3711_0[4:4], simp3711_0[5:5]);
  C3 I401 (simp3712_0[2:2], simp3711_0[6:6], simp3711_0[7:7], simp3711_0[8:8]);
  C2 I402 (simp3712_0[3:3], simp3711_0[9:9], simp3711_0[10:10]);
  C3 I403 (simp3713_0[0:0], simp3712_0[0:0], simp3712_0[1:1], simp3712_0[2:2]);
  BUFF I404 (simp3713_0[1:1], simp3712_0[3:3]);
  C2 I405 (icomp_2, simp3713_0[0:0], simp3713_0[1:1]);
  C2R I406 (choice_0, icomp_0, nchosen_0, reset);
  C2R I407 (choice_1, icomp_1, nchosen_0, reset);
  C2R I408 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I409 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I410 (nchosen_0, anychoice_0, o_0a);
  C2R I411 (i_0a, choice_0, o_0a, reset);
  C2R I412 (i_1a, choice_1, o_0a, reset);
  C2R I413 (i_2a, choice_2, o_0a, reset);
endmodule

// tkvr332_wo0w32_ro0w32o0w32o0w32o31w1 TeakV "r3" 32 [] [0] [0,0,0,31] [Many [32],Many [0],Many [0,0,0
//   ,0],Many [32,32,32,1]]
module tkvr332_wo0w32_ro0w32o0w32o0w32o31w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6021_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0, df_0[31:31], rg_3r);
  AND2 I521 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I522 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I523 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I524 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I525 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I526 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I527 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I528 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I529 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I530 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I531 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I532 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I533 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I534 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I535 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I536 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I537 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I538 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I539 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I540 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I541 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I542 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I543 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I544 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I545 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I546 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I547 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I548 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I549 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I550 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I551 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I552 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I553 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I554 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I555 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I556 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I557 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I558 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I559 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I560 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I561 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I562 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I563 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I564 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I565 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I566 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I567 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I568 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I569 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I570 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I571 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I572 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I573 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I574 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I575 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I576 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I577 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I578 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I579 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I580 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I581 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I582 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I583 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I584 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I585 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I586 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I587 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I588 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I589 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I590 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I591 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I592 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I593 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I594 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I595 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I596 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I597 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I598 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I599 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I600 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I601 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I602 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I603 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I604 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I605 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I606 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I607 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I608 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I609 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I610 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I611 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I612 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I613 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I614 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I615 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I616 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I617 (rd_3r1, dt_0[31:31], rg_3r);
  NOR3 I618 (simp6021_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I619 (simp6021_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I620 (simp6021_0[2:2], rg_2a, rg_3a);
  NAND3 I621 (anyread_0, simp6021_0[0:0], simp6021_0[1:1], simp6021_0[2:2]);
  BUFF I622 (wg_0a, wd_0a);
  BUFF I623 (rg_0a, rd_0a);
  BUFF I624 (rg_1a, rd_1a);
  BUFF I625 (rg_2a, rd_2a);
  BUFF I626 (rg_3a, rd_3a);
endmodule

// tkf32mo0w0_o0w32 TeakF [0,0] [One 32,Many [0,32]]
module tkf32mo0w0_o0w32 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I10 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I11 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I12 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I13 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I14 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I15 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I16 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I17 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I18 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I19 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I20 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I21 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I22 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I23 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I24 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I25 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I26 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I27 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I28 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I29 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I30 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I31 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I32 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I33 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I34 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I35 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I36 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I37 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I38 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I39 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I40 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I41 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I42 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I43 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I44 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I45 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I46 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I47 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I48 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I49 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I50 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I51 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I52 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I53 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I54 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I55 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I56 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I57 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I58 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I59 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I60 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I61 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I62 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I63 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I64 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I65 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I66 (o_0r, icomplete_0);
  C3 I67 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm2x32b TeakM [Many [32,32],One 32]
module tkm2x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2351_0;
  wire [3:0] simp2352_0;
  wire [1:0] simp2353_0;
  wire [31:0] comp1_0;
  wire [10:0] simp2691_0;
  wire [3:0] simp2692_0;
  wire [1:0] simp2693_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3]);
  OR2 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4]);
  OR2 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5]);
  OR2 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6]);
  OR2 I7 (o_0r0[7:7], gfint_0[7:7], gfint_1[7:7]);
  OR2 I8 (o_0r0[8:8], gfint_0[8:8], gfint_1[8:8]);
  OR2 I9 (o_0r0[9:9], gfint_0[9:9], gfint_1[9:9]);
  OR2 I10 (o_0r0[10:10], gfint_0[10:10], gfint_1[10:10]);
  OR2 I11 (o_0r0[11:11], gfint_0[11:11], gfint_1[11:11]);
  OR2 I12 (o_0r0[12:12], gfint_0[12:12], gfint_1[12:12]);
  OR2 I13 (o_0r0[13:13], gfint_0[13:13], gfint_1[13:13]);
  OR2 I14 (o_0r0[14:14], gfint_0[14:14], gfint_1[14:14]);
  OR2 I15 (o_0r0[15:15], gfint_0[15:15], gfint_1[15:15]);
  OR2 I16 (o_0r0[16:16], gfint_0[16:16], gfint_1[16:16]);
  OR2 I17 (o_0r0[17:17], gfint_0[17:17], gfint_1[17:17]);
  OR2 I18 (o_0r0[18:18], gfint_0[18:18], gfint_1[18:18]);
  OR2 I19 (o_0r0[19:19], gfint_0[19:19], gfint_1[19:19]);
  OR2 I20 (o_0r0[20:20], gfint_0[20:20], gfint_1[20:20]);
  OR2 I21 (o_0r0[21:21], gfint_0[21:21], gfint_1[21:21]);
  OR2 I22 (o_0r0[22:22], gfint_0[22:22], gfint_1[22:22]);
  OR2 I23 (o_0r0[23:23], gfint_0[23:23], gfint_1[23:23]);
  OR2 I24 (o_0r0[24:24], gfint_0[24:24], gfint_1[24:24]);
  OR2 I25 (o_0r0[25:25], gfint_0[25:25], gfint_1[25:25]);
  OR2 I26 (o_0r0[26:26], gfint_0[26:26], gfint_1[26:26]);
  OR2 I27 (o_0r0[27:27], gfint_0[27:27], gfint_1[27:27]);
  OR2 I28 (o_0r0[28:28], gfint_0[28:28], gfint_1[28:28]);
  OR2 I29 (o_0r0[29:29], gfint_0[29:29], gfint_1[29:29]);
  OR2 I30 (o_0r0[30:30], gfint_0[30:30], gfint_1[30:30]);
  OR2 I31 (o_0r0[31:31], gfint_0[31:31], gfint_1[31:31]);
  OR2 I32 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I33 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I34 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  OR2 I35 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3]);
  OR2 I36 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4]);
  OR2 I37 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5]);
  OR2 I38 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6]);
  OR2 I39 (o_0r1[7:7], gtint_0[7:7], gtint_1[7:7]);
  OR2 I40 (o_0r1[8:8], gtint_0[8:8], gtint_1[8:8]);
  OR2 I41 (o_0r1[9:9], gtint_0[9:9], gtint_1[9:9]);
  OR2 I42 (o_0r1[10:10], gtint_0[10:10], gtint_1[10:10]);
  OR2 I43 (o_0r1[11:11], gtint_0[11:11], gtint_1[11:11]);
  OR2 I44 (o_0r1[12:12], gtint_0[12:12], gtint_1[12:12]);
  OR2 I45 (o_0r1[13:13], gtint_0[13:13], gtint_1[13:13]);
  OR2 I46 (o_0r1[14:14], gtint_0[14:14], gtint_1[14:14]);
  OR2 I47 (o_0r1[15:15], gtint_0[15:15], gtint_1[15:15]);
  OR2 I48 (o_0r1[16:16], gtint_0[16:16], gtint_1[16:16]);
  OR2 I49 (o_0r1[17:17], gtint_0[17:17], gtint_1[17:17]);
  OR2 I50 (o_0r1[18:18], gtint_0[18:18], gtint_1[18:18]);
  OR2 I51 (o_0r1[19:19], gtint_0[19:19], gtint_1[19:19]);
  OR2 I52 (o_0r1[20:20], gtint_0[20:20], gtint_1[20:20]);
  OR2 I53 (o_0r1[21:21], gtint_0[21:21], gtint_1[21:21]);
  OR2 I54 (o_0r1[22:22], gtint_0[22:22], gtint_1[22:22]);
  OR2 I55 (o_0r1[23:23], gtint_0[23:23], gtint_1[23:23]);
  OR2 I56 (o_0r1[24:24], gtint_0[24:24], gtint_1[24:24]);
  OR2 I57 (o_0r1[25:25], gtint_0[25:25], gtint_1[25:25]);
  OR2 I58 (o_0r1[26:26], gtint_0[26:26], gtint_1[26:26]);
  OR2 I59 (o_0r1[27:27], gtint_0[27:27], gtint_1[27:27]);
  OR2 I60 (o_0r1[28:28], gtint_0[28:28], gtint_1[28:28]);
  OR2 I61 (o_0r1[29:29], gtint_0[29:29], gtint_1[29:29]);
  OR2 I62 (o_0r1[30:30], gtint_0[30:30], gtint_1[30:30]);
  OR2 I63 (o_0r1[31:31], gtint_0[31:31], gtint_1[31:31]);
  AND2 I64 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I65 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I66 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I67 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I68 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I69 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I70 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I71 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I72 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I73 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I74 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I75 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I76 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I77 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I78 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I79 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I80 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I81 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I82 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I83 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I84 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I85 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I86 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I87 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I88 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I89 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I90 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I91 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I92 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I93 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I94 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I95 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I96 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I97 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I98 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I99 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I100 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I101 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I102 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I103 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I104 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I105 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I106 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I107 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I108 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I109 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I110 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I111 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I112 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I113 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I114 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I115 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I116 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I117 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I118 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I119 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I120 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I121 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I122 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I123 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I124 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I125 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I126 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I127 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I128 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I129 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I130 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I131 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I132 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I133 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I134 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I135 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I136 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I137 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I138 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I139 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I140 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I141 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I142 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I143 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I144 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I145 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I146 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I147 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I148 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I149 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I150 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I151 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I152 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I153 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I154 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I155 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I156 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I157 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I158 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I159 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I160 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I161 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I162 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I163 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I164 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I165 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I166 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I167 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I168 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I169 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I170 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I171 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I172 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I173 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I174 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I175 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I176 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I177 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I178 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I179 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I180 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I181 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I182 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I183 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I184 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I185 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I186 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I187 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I188 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I189 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I190 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I191 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  OR2 I192 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I193 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I194 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I195 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I196 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I197 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I198 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I199 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I200 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I201 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I202 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I203 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I204 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I205 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I206 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I207 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I208 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I209 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I210 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I211 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I212 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I213 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I214 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I215 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I216 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I217 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I218 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I219 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I220 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I221 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I222 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I223 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I224 (simp2351_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I225 (simp2351_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I226 (simp2351_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I227 (simp2351_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I228 (simp2351_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I229 (simp2351_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I230 (simp2351_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I231 (simp2351_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I232 (simp2351_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I233 (simp2351_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I234 (simp2351_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I235 (simp2352_0[0:0], simp2351_0[0:0], simp2351_0[1:1], simp2351_0[2:2]);
  C3 I236 (simp2352_0[1:1], simp2351_0[3:3], simp2351_0[4:4], simp2351_0[5:5]);
  C3 I237 (simp2352_0[2:2], simp2351_0[6:6], simp2351_0[7:7], simp2351_0[8:8]);
  C2 I238 (simp2352_0[3:3], simp2351_0[9:9], simp2351_0[10:10]);
  C3 I239 (simp2353_0[0:0], simp2352_0[0:0], simp2352_0[1:1], simp2352_0[2:2]);
  BUFF I240 (simp2353_0[1:1], simp2352_0[3:3]);
  C2 I241 (icomp_0, simp2353_0[0:0], simp2353_0[1:1]);
  OR2 I242 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I243 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I244 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I245 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I246 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I247 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I248 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I249 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I250 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I251 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I252 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I253 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I254 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I255 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I256 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I257 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I258 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I259 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I260 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I261 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I262 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I263 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I264 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I265 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I266 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I267 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I268 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I269 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I270 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I271 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I272 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I273 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I274 (simp2691_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I275 (simp2691_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I276 (simp2691_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I277 (simp2691_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I278 (simp2691_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I279 (simp2691_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I280 (simp2691_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I281 (simp2691_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I282 (simp2691_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I283 (simp2691_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I284 (simp2691_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I285 (simp2692_0[0:0], simp2691_0[0:0], simp2691_0[1:1], simp2691_0[2:2]);
  C3 I286 (simp2692_0[1:1], simp2691_0[3:3], simp2691_0[4:4], simp2691_0[5:5]);
  C3 I287 (simp2692_0[2:2], simp2691_0[6:6], simp2691_0[7:7], simp2691_0[8:8]);
  C2 I288 (simp2692_0[3:3], simp2691_0[9:9], simp2691_0[10:10]);
  C3 I289 (simp2693_0[0:0], simp2692_0[0:0], simp2692_0[1:1], simp2692_0[2:2]);
  BUFF I290 (simp2693_0[1:1], simp2692_0[3:3]);
  C2 I291 (icomp_1, simp2693_0[0:0], simp2693_0[1:1]);
  C2R I292 (choice_0, icomp_0, nchosen_0, reset);
  C2R I293 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I294 (anychoice_0, choice_0, choice_1);
  NOR2 I295 (nchosen_0, anychoice_0, o_0a);
  C2R I296 (i_0a, choice_0, o_0a, reset);
  C2R I297 (i_1a, choice_1, o_0a, reset);
endmodule

// tko0m2_1nm2b1 TeakO [
//     (1,TeakOConstant 2 1)] [One 0,One 2]
module tko0m2_1nm2b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  GND I3 (o_0r1[1:1]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tko0m2_1nm2b2 TeakO [
//     (1,TeakOConstant 2 2)] [One 0,One 2]
module tko0m2_1nm2b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  GND I3 (o_0r1[0:0]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tkm2x2b TeakM [Many [2,2],One 2]
module tkm2x2b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire [1:0] gfint_0;
  wire [1:0] gfint_1;
  wire [1:0] gtint_0;
  wire [1:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [1:0] comp0_0;
  wire [1:0] comp1_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I3 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  AND2 I4 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I5 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I6 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I7 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I8 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I9 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I10 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I11 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  OR2 I12 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I13 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I14 (icomp_0, comp0_0[0:0], comp0_0[1:1]);
  OR2 I15 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I16 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  C2 I17 (icomp_1, comp1_0[0:0], comp1_0[1:1]);
  C2R I18 (choice_0, icomp_0, nchosen_0, reset);
  C2R I19 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I20 (anychoice_0, choice_0, choice_1);
  NOR2 I21 (nchosen_0, anychoice_0, o_0a);
  C2R I22 (i_0a, choice_0, o_0a, reset);
  C2R I23 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj2m0_2 TeakJ [Many [0,2],One 2]
module tkj2m0_2 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [1:0] joinf_0;
  wire [1:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joint_0[0:0], i_1r1[0:0]);
  BUFF I3 (joint_0[1:1], i_1r1[1:1]);
  BUFF I4 (icomplete_0, i_0r);
  C2 I5 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I6 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I7 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I8 (o_0r1[1:1], joint_0[1:1]);
  BUFF I9 (i_0a, o_0a);
  BUFF I10 (i_1a, o_0a);
endmodule

// tks2_o0w2_1o0w0_2o0w0 TeakS (0+:2) [([Imp 1 0],0),([Imp 2 0],0)] [One 2,Many [0,0]]
module tks2_o0w2_1o0w0_2o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire [1:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[0:0], i_0r0[1:1]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r0[0:0], i_0r1[1:1]);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I7 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I8 (icomplete_0, comp_0[0:0], comp_0[1:1]);
  BUFF I9 (o_0r, gsel_0);
  BUFF I10 (o_1r, gsel_1);
  OR2 I11 (oack_0, o_0a, o_1a);
  C2 I12 (i_0a, oack_0, icomplete_0);
endmodule

// tkvr232_wo0w32_ro0w32o0w32o31w1 TeakV "r2" 32 [] [0] [0,0,31] [Many [32],Many [0],Many [0,0,0],Many 
//   [32,32,1]]
module tkvr232_wo0w32_ro0w32o0w32o31w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp5381_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0, df_0[31:31], rg_2r);
  AND2 I489 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I490 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I491 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I492 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I493 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I494 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I495 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I496 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I497 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I498 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I499 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I500 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I501 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I502 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I503 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I504 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I505 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I506 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I507 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I508 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I509 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I510 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I511 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I512 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I513 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I514 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I515 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I516 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I517 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I518 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I519 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I520 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I521 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I522 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I523 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I524 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I525 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I526 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I527 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I528 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I529 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I530 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I531 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I532 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I533 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I534 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I535 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I536 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I537 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I538 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I539 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I540 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I541 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I542 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I543 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I544 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I545 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I546 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I547 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I548 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I549 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I550 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I551 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I552 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I553 (rd_2r1, dt_0[31:31], rg_2r);
  NOR3 I554 (simp5381_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I555 (simp5381_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I556 (anyread_0, simp5381_0[0:0], simp5381_0[1:1]);
  BUFF I557 (wg_0a, wd_0a);
  BUFF I558 (rg_0a, rd_0a);
  BUFF I559 (rg_1a, rd_1a);
  BUFF I560 (rg_2a, rd_2a);
endmodule

// tkvr132_wo0w32_ro0w32o0w32o0w32 TeakV "r1" 32 [] [0] [0,0,0] [Many [32],Many [0],Many [0,0,0],Many [
//   32,32,32]]
module tkvr132_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tks32_o0w32_3cfffffffcm4cfffffff8m5cfffffff8m6cfffffff8m8cfffffff0m9cfffffff0macfffffff0m10cffffffe0
//   m11cffffffe0m12cffffffe0m20cffffffc0m21cffffffc0m22cffffffc0m40cffffff80m41cffffff80m42cffffff80m80c
//   ffffff00m81cffffff00m82cffffff00m100cfffffe00m101cfffffe00m102cfffffe00m200cfffffc00m201cfffffc00m20
//   2cfffffc00m400cfffff800m401cfffff800m402cfffff800m800cfffff000m801cfffff000m802cfffff000m1000cffffe0
//   00m1001cffffe000m1002cffffe000m2000cffffc000m2001cffffc000m2002cffffc000m4000cffff8000m4001cffff8000
//   m4002cffff8000m8000cffff0000m8001cffff0000m8002cffff0000m10000cfffe0000m10001cfffe0000m10002cfffe000
//   0m20000cfffc0000m20001cfffc0000m20002cfffc0000m40000cfff80000m40001cfff80000m40002cfff80000m80000cff
//   f00000m80001cfff00000m80002cfff00000m100000cffe00000m100001cffe00000m100002cffe00000m200000cffc00000
//   m200001cffc00000m200002cffc00000m400000cff800000m400001cff800000m400002cff800000m800000cff000000m800
//   001cff000000m800002cff000000m1000000cfe000000m1000001cfe000000m1000002cfe000000m2000000cfc000000m200
//   0001cfc000000m2000002cfc000000m4000000cf8000000m4000001cf8000000m4000002cf8000000m8000000cf0000000m8
//   000001cf0000000m8000002cf0000000m10000000ce0000000m10000001ce0000000m10000002ce0000000m20000000cc000
//   0000m20000001cc0000000m20000002cc0000000m40000000c80000000m40000001c80000000m40000002c80000000m80000
//   000m80000001m80000002o0w0_0o0w0_1o0w0_2o0w0 TeakS (0+:32) [([Imp 3 4294967292,Imp 4 4294967288,Imp 5
//    4294967288,Imp 6 4294967288,Imp 8 4294967280,Imp 9 4294967280,Imp 10 4294967280,Imp 16 4294967264,I
//   mp 17 4294967264,Imp 18 4294967264,Imp 32 4294967232,Imp 33 4294967232,Imp 34 4294967232,Imp 64 4294
//   967168,Imp 65 4294967168,Imp 66 4294967168,Imp 128 4294967040,Imp 129 4294967040,Imp 130 4294967040,
//   Imp 256 4294966784,Imp 257 4294966784,Imp 258 4294966784,Imp 512 4294966272,Imp 513 4294966272,Imp 5
//   14 4294966272,Imp 1024 4294965248,Imp 1025 4294965248,Imp 1026 4294965248,Imp 2048 4294963200,Imp 20
//   49 4294963200,Imp 2050 4294963200,Imp 4096 4294959104,Imp 4097 4294959104,Imp 4098 4294959104,Imp 81
//   92 4294950912,Imp 8193 4294950912,Imp 8194 4294950912,Imp 16384 4294934528,Imp 16385 4294934528,Imp 
//   16386 4294934528,Imp 32768 4294901760,Imp 32769 4294901760,Imp 32770 4294901760,Imp 65536 4294836224
//   ,Imp 65537 4294836224,Imp 65538 4294836224,Imp 131072 4294705152,Imp 131073 4294705152,Imp 131074 42
//   94705152,Imp 262144 4294443008,Imp 262145 4294443008,Imp 262146 4294443008,Imp 524288 4293918720,Imp
//    524289 4293918720,Imp 524290 4293918720,Imp 1048576 4292870144,Imp 1048577 4292870144,Imp 1048578 4
//   292870144,Imp 2097152 4290772992,Imp 2097153 4290772992,Imp 2097154 4290772992,Imp 4194304 428657868
//   8,Imp 4194305 4286578688,Imp 4194306 4286578688,Imp 8388608 4278190080,Imp 8388609 4278190080,Imp 83
//   88610 4278190080,Imp 16777216 4261412864,Imp 16777217 4261412864,Imp 16777218 4261412864,Imp 3355443
//   2 4227858432,Imp 33554433 4227858432,Imp 33554434 4227858432,Imp 67108864 4160749568,Imp 67108865 41
//   60749568,Imp 67108866 4160749568,Imp 134217728 4026531840,Imp 134217729 4026531840,Imp 134217730 402
//   6531840,Imp 268435456 3758096384,Imp 268435457 3758096384,Imp 268435458 3758096384,Imp 536870912 322
//   1225472,Imp 536870913 3221225472,Imp 536870914 3221225472,Imp 1073741824 2147483648,Imp 1073741825 2
//   147483648,Imp 1073741826 2147483648,Imp 2147483648 0,Imp 2147483649 0,Imp 2147483650 0],0),([Imp 0 0
//   ],0),([Imp 1 0],0),([Imp 2 0],0)] [One 32,Many [0,0,0,0]]
module tks32_o0w32_3cfffffffcm4cfffffff8m5cfffffff8m6cfffffff8m8cfffffff0m9cfffffff0macfffffff0m10cffffffe0m11cffffffe0m12cffffffe0m20cffffffc0m21cffffffc0m22cffffffc0m40cffffff80m41cffffff80m42cffffff80m80cffffff00m81cffffff00m82cffffff00m100cfffffe00m101cfffffe00m102cfffffe00m200cfffffc00m201cfffffc00m202cfffffc00m400cfffff800m401cfffff800m402cfffff800m800cfffff000m801cfffff000m802cfffff000m1000cffffe000m1001cffffe000m1002cffffe000m2000cffffc000m2001cffffc000m2002cffffc000m4000cffff8000m4001cffff8000m4002cffff8000m8000cffff0000m8001cffff0000m8002cffff0000m10000cfffe0000m10001cfffe0000m10002cfffe0000m20000cfffc0000m20001cfffc0000m20002cfffc0000m40000cfff80000m40001cfff80000m40002cfff80000m80000cfff00000m80001cfff00000m80002cfff00000m100000cffe00000m100001cffe00000m100002cffe00000m200000cffc00000m200001cffc00000m200002cffc00000m400000cff800000m400001cff800000m400002cff800000m800000cff000000m800001cff000000m800002cff000000m1000000cfe000000m1000001cfe000000m1000002cfe000000m2000000cfc000000m2000001cfc000000m2000002cfc000000m4000000cf8000000m4000001cf8000000m4000002cf8000000m8000000cf0000000m8000001cf0000000m8000002cf0000000m10000000ce0000000m10000001ce0000000m10000002ce0000000m20000000cc0000000m20000001cc0000000m20000002cc0000000m40000000c80000000m40000001c80000000m40000002c80000000m80000000m80000001m80000002o0w0_0o0w0_1o0w0_2o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire oack_0;
  wire [90:0] match0_0;
  wire [30:0] simp111_0;
  wire [10:0] simp112_0;
  wire [3:0] simp113_0;
  wire [1:0] simp114_0;
  wire [1:0] simp161_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [2:0] simp251_0;
  wire [2:0] simp261_0;
  wire [2:0] simp271_0;
  wire [2:0] simp281_0;
  wire [2:0] simp291_0;
  wire [2:0] simp301_0;
  wire [2:0] simp311_0;
  wire [2:0] simp321_0;
  wire [2:0] simp331_0;
  wire [3:0] simp341_0;
  wire [1:0] simp342_0;
  wire [3:0] simp351_0;
  wire [1:0] simp352_0;
  wire [3:0] simp361_0;
  wire [1:0] simp362_0;
  wire [3:0] simp371_0;
  wire [1:0] simp372_0;
  wire [3:0] simp381_0;
  wire [1:0] simp382_0;
  wire [3:0] simp391_0;
  wire [1:0] simp392_0;
  wire [3:0] simp401_0;
  wire [1:0] simp402_0;
  wire [3:0] simp411_0;
  wire [1:0] simp412_0;
  wire [3:0] simp421_0;
  wire [1:0] simp422_0;
  wire [4:0] simp431_0;
  wire [1:0] simp432_0;
  wire [4:0] simp441_0;
  wire [1:0] simp442_0;
  wire [4:0] simp451_0;
  wire [1:0] simp452_0;
  wire [4:0] simp461_0;
  wire [1:0] simp462_0;
  wire [4:0] simp471_0;
  wire [1:0] simp472_0;
  wire [4:0] simp481_0;
  wire [1:0] simp482_0;
  wire [4:0] simp491_0;
  wire [1:0] simp492_0;
  wire [4:0] simp501_0;
  wire [1:0] simp502_0;
  wire [4:0] simp511_0;
  wire [1:0] simp512_0;
  wire [5:0] simp521_0;
  wire [1:0] simp522_0;
  wire [5:0] simp531_0;
  wire [1:0] simp532_0;
  wire [5:0] simp541_0;
  wire [1:0] simp542_0;
  wire [5:0] simp551_0;
  wire [1:0] simp552_0;
  wire [5:0] simp561_0;
  wire [1:0] simp562_0;
  wire [5:0] simp571_0;
  wire [1:0] simp572_0;
  wire [5:0] simp581_0;
  wire [1:0] simp582_0;
  wire [5:0] simp591_0;
  wire [1:0] simp592_0;
  wire [5:0] simp601_0;
  wire [1:0] simp602_0;
  wire [6:0] simp611_0;
  wire [2:0] simp612_0;
  wire [6:0] simp621_0;
  wire [2:0] simp622_0;
  wire [6:0] simp631_0;
  wire [2:0] simp632_0;
  wire [6:0] simp641_0;
  wire [2:0] simp642_0;
  wire [6:0] simp651_0;
  wire [2:0] simp652_0;
  wire [6:0] simp661_0;
  wire [2:0] simp662_0;
  wire [6:0] simp671_0;
  wire [2:0] simp672_0;
  wire [6:0] simp681_0;
  wire [2:0] simp682_0;
  wire [6:0] simp691_0;
  wire [2:0] simp692_0;
  wire [7:0] simp701_0;
  wire [2:0] simp702_0;
  wire [7:0] simp711_0;
  wire [2:0] simp712_0;
  wire [7:0] simp721_0;
  wire [2:0] simp722_0;
  wire [7:0] simp731_0;
  wire [2:0] simp732_0;
  wire [7:0] simp741_0;
  wire [2:0] simp742_0;
  wire [7:0] simp751_0;
  wire [2:0] simp752_0;
  wire [7:0] simp761_0;
  wire [2:0] simp762_0;
  wire [7:0] simp771_0;
  wire [2:0] simp772_0;
  wire [7:0] simp781_0;
  wire [2:0] simp782_0;
  wire [8:0] simp791_0;
  wire [2:0] simp792_0;
  wire [8:0] simp801_0;
  wire [2:0] simp802_0;
  wire [8:0] simp811_0;
  wire [2:0] simp812_0;
  wire [8:0] simp821_0;
  wire [2:0] simp822_0;
  wire [8:0] simp831_0;
  wire [2:0] simp832_0;
  wire [8:0] simp841_0;
  wire [2:0] simp842_0;
  wire [8:0] simp851_0;
  wire [2:0] simp852_0;
  wire [8:0] simp861_0;
  wire [2:0] simp862_0;
  wire [8:0] simp871_0;
  wire [2:0] simp872_0;
  wire [9:0] simp881_0;
  wire [3:0] simp882_0;
  wire [1:0] simp883_0;
  wire [9:0] simp891_0;
  wire [3:0] simp892_0;
  wire [1:0] simp893_0;
  wire [9:0] simp901_0;
  wire [3:0] simp902_0;
  wire [1:0] simp903_0;
  wire [9:0] simp911_0;
  wire [3:0] simp912_0;
  wire [1:0] simp913_0;
  wire [9:0] simp921_0;
  wire [3:0] simp922_0;
  wire [1:0] simp923_0;
  wire [9:0] simp931_0;
  wire [3:0] simp932_0;
  wire [1:0] simp933_0;
  wire [9:0] simp941_0;
  wire [3:0] simp942_0;
  wire [1:0] simp943_0;
  wire [9:0] simp951_0;
  wire [3:0] simp952_0;
  wire [1:0] simp953_0;
  wire [9:0] simp961_0;
  wire [3:0] simp962_0;
  wire [1:0] simp963_0;
  wire [10:0] simp971_0;
  wire [3:0] simp972_0;
  wire [1:0] simp973_0;
  wire [10:0] simp981_0;
  wire [3:0] simp982_0;
  wire [1:0] simp983_0;
  wire [10:0] simp991_0;
  wire [3:0] simp992_0;
  wire [1:0] simp993_0;
  wire [10:0] simp1001_0;
  wire [3:0] simp1002_0;
  wire [1:0] simp1003_0;
  wire [10:0] simp1011_0;
  wire [3:0] simp1012_0;
  wire [1:0] simp1013_0;
  wire [10:0] simp1021_0;
  wire [3:0] simp1022_0;
  wire [1:0] simp1023_0;
  wire match1_0;
  wire [10:0] simp1051_0;
  wire [3:0] simp1052_0;
  wire [1:0] simp1053_0;
  wire match2_0;
  wire [10:0] simp1081_0;
  wire [3:0] simp1082_0;
  wire [1:0] simp1083_0;
  wire match3_0;
  wire [10:0] simp1111_0;
  wire [3:0] simp1112_0;
  wire [1:0] simp1113_0;
  wire [31:0] comp_0;
  wire [10:0] simp1491_0;
  wire [3:0] simp1492_0;
  wire [1:0] simp1493_0;
  wire [1:0] simp1541_0;
  NOR3 I0 (simp111_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp111_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NOR3 I2 (simp111_0[2:2], match0_0[6:6], match0_0[7:7], match0_0[8:8]);
  NOR3 I3 (simp111_0[3:3], match0_0[9:9], match0_0[10:10], match0_0[11:11]);
  NOR3 I4 (simp111_0[4:4], match0_0[12:12], match0_0[13:13], match0_0[14:14]);
  NOR3 I5 (simp111_0[5:5], match0_0[15:15], match0_0[16:16], match0_0[17:17]);
  NOR3 I6 (simp111_0[6:6], match0_0[18:18], match0_0[19:19], match0_0[20:20]);
  NOR3 I7 (simp111_0[7:7], match0_0[21:21], match0_0[22:22], match0_0[23:23]);
  NOR3 I8 (simp111_0[8:8], match0_0[24:24], match0_0[25:25], match0_0[26:26]);
  NOR3 I9 (simp111_0[9:9], match0_0[27:27], match0_0[28:28], match0_0[29:29]);
  NOR3 I10 (simp111_0[10:10], match0_0[30:30], match0_0[31:31], match0_0[32:32]);
  NOR3 I11 (simp111_0[11:11], match0_0[33:33], match0_0[34:34], match0_0[35:35]);
  NOR3 I12 (simp111_0[12:12], match0_0[36:36], match0_0[37:37], match0_0[38:38]);
  NOR3 I13 (simp111_0[13:13], match0_0[39:39], match0_0[40:40], match0_0[41:41]);
  NOR3 I14 (simp111_0[14:14], match0_0[42:42], match0_0[43:43], match0_0[44:44]);
  NOR3 I15 (simp111_0[15:15], match0_0[45:45], match0_0[46:46], match0_0[47:47]);
  NOR3 I16 (simp111_0[16:16], match0_0[48:48], match0_0[49:49], match0_0[50:50]);
  NOR3 I17 (simp111_0[17:17], match0_0[51:51], match0_0[52:52], match0_0[53:53]);
  NOR3 I18 (simp111_0[18:18], match0_0[54:54], match0_0[55:55], match0_0[56:56]);
  NOR3 I19 (simp111_0[19:19], match0_0[57:57], match0_0[58:58], match0_0[59:59]);
  NOR3 I20 (simp111_0[20:20], match0_0[60:60], match0_0[61:61], match0_0[62:62]);
  NOR3 I21 (simp111_0[21:21], match0_0[63:63], match0_0[64:64], match0_0[65:65]);
  NOR3 I22 (simp111_0[22:22], match0_0[66:66], match0_0[67:67], match0_0[68:68]);
  NOR3 I23 (simp111_0[23:23], match0_0[69:69], match0_0[70:70], match0_0[71:71]);
  NOR3 I24 (simp111_0[24:24], match0_0[72:72], match0_0[73:73], match0_0[74:74]);
  NOR3 I25 (simp111_0[25:25], match0_0[75:75], match0_0[76:76], match0_0[77:77]);
  NOR3 I26 (simp111_0[26:26], match0_0[78:78], match0_0[79:79], match0_0[80:80]);
  NOR3 I27 (simp111_0[27:27], match0_0[81:81], match0_0[82:82], match0_0[83:83]);
  NOR3 I28 (simp111_0[28:28], match0_0[84:84], match0_0[85:85], match0_0[86:86]);
  NOR3 I29 (simp111_0[29:29], match0_0[87:87], match0_0[88:88], match0_0[89:89]);
  INV I30 (simp111_0[30:30], match0_0[90:90]);
  NAND3 I31 (simp112_0[0:0], simp111_0[0:0], simp111_0[1:1], simp111_0[2:2]);
  NAND3 I32 (simp112_0[1:1], simp111_0[3:3], simp111_0[4:4], simp111_0[5:5]);
  NAND3 I33 (simp112_0[2:2], simp111_0[6:6], simp111_0[7:7], simp111_0[8:8]);
  NAND3 I34 (simp112_0[3:3], simp111_0[9:9], simp111_0[10:10], simp111_0[11:11]);
  NAND3 I35 (simp112_0[4:4], simp111_0[12:12], simp111_0[13:13], simp111_0[14:14]);
  NAND3 I36 (simp112_0[5:5], simp111_0[15:15], simp111_0[16:16], simp111_0[17:17]);
  NAND3 I37 (simp112_0[6:6], simp111_0[18:18], simp111_0[19:19], simp111_0[20:20]);
  NAND3 I38 (simp112_0[7:7], simp111_0[21:21], simp111_0[22:22], simp111_0[23:23]);
  NAND3 I39 (simp112_0[8:8], simp111_0[24:24], simp111_0[25:25], simp111_0[26:26]);
  NAND3 I40 (simp112_0[9:9], simp111_0[27:27], simp111_0[28:28], simp111_0[29:29]);
  INV I41 (simp112_0[10:10], simp111_0[30:30]);
  NOR3 I42 (simp113_0[0:0], simp112_0[0:0], simp112_0[1:1], simp112_0[2:2]);
  NOR3 I43 (simp113_0[1:1], simp112_0[3:3], simp112_0[4:4], simp112_0[5:5]);
  NOR3 I44 (simp113_0[2:2], simp112_0[6:6], simp112_0[7:7], simp112_0[8:8]);
  NOR2 I45 (simp113_0[3:3], simp112_0[9:9], simp112_0[10:10]);
  NAND3 I46 (simp114_0[0:0], simp113_0[0:0], simp113_0[1:1], simp113_0[2:2]);
  INV I47 (simp114_0[1:1], simp113_0[3:3]);
  OR2 I48 (sel_0, simp114_0[0:0], simp114_0[1:1]);
  C2 I49 (match0_0[0:0], i_0r1[0:0], i_0r1[1:1]);
  C3 I50 (match0_0[1:1], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I51 (match0_0[2:2], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I52 (match0_0[3:3], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I53 (simp161_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I54 (simp161_0[1:1], i_0r1[3:3]);
  C2 I55 (match0_0[4:4], simp161_0[0:0], simp161_0[1:1]);
  C3 I56 (simp171_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I57 (simp171_0[1:1], i_0r1[3:3]);
  C2 I58 (match0_0[5:5], simp171_0[0:0], simp171_0[1:1]);
  C3 I59 (simp181_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I60 (simp181_0[1:1], i_0r1[3:3]);
  C2 I61 (match0_0[6:6], simp181_0[0:0], simp181_0[1:1]);
  C3 I62 (simp191_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I63 (simp191_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I64 (match0_0[7:7], simp191_0[0:0], simp191_0[1:1]);
  C3 I65 (simp201_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I66 (simp201_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I67 (match0_0[8:8], simp201_0[0:0], simp201_0[1:1]);
  C3 I68 (simp211_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C2 I69 (simp211_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I70 (match0_0[9:9], simp211_0[0:0], simp211_0[1:1]);
  C3 I71 (simp221_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I72 (simp221_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I73 (match0_0[10:10], simp221_0[0:0], simp221_0[1:1]);
  C3 I74 (simp231_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I75 (simp231_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I76 (match0_0[11:11], simp231_0[0:0], simp231_0[1:1]);
  C3 I77 (simp241_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I78 (simp241_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I79 (match0_0[12:12], simp241_0[0:0], simp241_0[1:1]);
  C3 I80 (simp251_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I81 (simp251_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I82 (simp251_0[2:2], i_0r1[6:6]);
  C3 I83 (match0_0[13:13], simp251_0[0:0], simp251_0[1:1], simp251_0[2:2]);
  C3 I84 (simp261_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I85 (simp261_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I86 (simp261_0[2:2], i_0r1[6:6]);
  C3 I87 (match0_0[14:14], simp261_0[0:0], simp261_0[1:1], simp261_0[2:2]);
  C3 I88 (simp271_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I89 (simp271_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I90 (simp271_0[2:2], i_0r1[6:6]);
  C3 I91 (match0_0[15:15], simp271_0[0:0], simp271_0[1:1], simp271_0[2:2]);
  C3 I92 (simp281_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I93 (simp281_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I94 (simp281_0[2:2], i_0r0[6:6], i_0r1[7:7]);
  C3 I95 (match0_0[16:16], simp281_0[0:0], simp281_0[1:1], simp281_0[2:2]);
  C3 I96 (simp291_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I97 (simp291_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I98 (simp291_0[2:2], i_0r0[6:6], i_0r1[7:7]);
  C3 I99 (match0_0[17:17], simp291_0[0:0], simp291_0[1:1], simp291_0[2:2]);
  C3 I100 (simp301_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I101 (simp301_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I102 (simp301_0[2:2], i_0r0[6:6], i_0r1[7:7]);
  C3 I103 (match0_0[18:18], simp301_0[0:0], simp301_0[1:1], simp301_0[2:2]);
  C3 I104 (simp311_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I105 (simp311_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I106 (simp311_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r1[8:8]);
  C3 I107 (match0_0[19:19], simp311_0[0:0], simp311_0[1:1], simp311_0[2:2]);
  C3 I108 (simp321_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I109 (simp321_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I110 (simp321_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r1[8:8]);
  C3 I111 (match0_0[20:20], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  C3 I112 (simp331_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I113 (simp331_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I114 (simp331_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r1[8:8]);
  C3 I115 (match0_0[21:21], simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  C3 I116 (simp341_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I117 (simp341_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I118 (simp341_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  BUFF I119 (simp341_0[3:3], i_0r1[9:9]);
  C3 I120 (simp342_0[0:0], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  BUFF I121 (simp342_0[1:1], simp341_0[3:3]);
  C2 I122 (match0_0[22:22], simp342_0[0:0], simp342_0[1:1]);
  C3 I123 (simp351_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I124 (simp351_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I125 (simp351_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  BUFF I126 (simp351_0[3:3], i_0r1[9:9]);
  C3 I127 (simp352_0[0:0], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  BUFF I128 (simp352_0[1:1], simp351_0[3:3]);
  C2 I129 (match0_0[23:23], simp352_0[0:0], simp352_0[1:1]);
  C3 I130 (simp361_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I131 (simp361_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I132 (simp361_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  BUFF I133 (simp361_0[3:3], i_0r1[9:9]);
  C3 I134 (simp362_0[0:0], simp361_0[0:0], simp361_0[1:1], simp361_0[2:2]);
  BUFF I135 (simp362_0[1:1], simp361_0[3:3]);
  C2 I136 (match0_0[24:24], simp362_0[0:0], simp362_0[1:1]);
  C3 I137 (simp371_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I138 (simp371_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I139 (simp371_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I140 (simp371_0[3:3], i_0r0[9:9], i_0r1[10:10]);
  C3 I141 (simp372_0[0:0], simp371_0[0:0], simp371_0[1:1], simp371_0[2:2]);
  BUFF I142 (simp372_0[1:1], simp371_0[3:3]);
  C2 I143 (match0_0[25:25], simp372_0[0:0], simp372_0[1:1]);
  C3 I144 (simp381_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I145 (simp381_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I146 (simp381_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I147 (simp381_0[3:3], i_0r0[9:9], i_0r1[10:10]);
  C3 I148 (simp382_0[0:0], simp381_0[0:0], simp381_0[1:1], simp381_0[2:2]);
  BUFF I149 (simp382_0[1:1], simp381_0[3:3]);
  C2 I150 (match0_0[26:26], simp382_0[0:0], simp382_0[1:1]);
  C3 I151 (simp391_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I152 (simp391_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I153 (simp391_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I154 (simp391_0[3:3], i_0r0[9:9], i_0r1[10:10]);
  C3 I155 (simp392_0[0:0], simp391_0[0:0], simp391_0[1:1], simp391_0[2:2]);
  BUFF I156 (simp392_0[1:1], simp391_0[3:3]);
  C2 I157 (match0_0[27:27], simp392_0[0:0], simp392_0[1:1]);
  C3 I158 (simp401_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I159 (simp401_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I160 (simp401_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I161 (simp401_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r1[11:11]);
  C3 I162 (simp402_0[0:0], simp401_0[0:0], simp401_0[1:1], simp401_0[2:2]);
  BUFF I163 (simp402_0[1:1], simp401_0[3:3]);
  C2 I164 (match0_0[28:28], simp402_0[0:0], simp402_0[1:1]);
  C3 I165 (simp411_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I166 (simp411_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I167 (simp411_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I168 (simp411_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r1[11:11]);
  C3 I169 (simp412_0[0:0], simp411_0[0:0], simp411_0[1:1], simp411_0[2:2]);
  BUFF I170 (simp412_0[1:1], simp411_0[3:3]);
  C2 I171 (match0_0[29:29], simp412_0[0:0], simp412_0[1:1]);
  C3 I172 (simp421_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I173 (simp421_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I174 (simp421_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I175 (simp421_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r1[11:11]);
  C3 I176 (simp422_0[0:0], simp421_0[0:0], simp421_0[1:1], simp421_0[2:2]);
  BUFF I177 (simp422_0[1:1], simp421_0[3:3]);
  C2 I178 (match0_0[30:30], simp422_0[0:0], simp422_0[1:1]);
  C3 I179 (simp431_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I180 (simp431_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I181 (simp431_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I182 (simp431_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  BUFF I183 (simp431_0[4:4], i_0r1[12:12]);
  C3 I184 (simp432_0[0:0], simp431_0[0:0], simp431_0[1:1], simp431_0[2:2]);
  C2 I185 (simp432_0[1:1], simp431_0[3:3], simp431_0[4:4]);
  C2 I186 (match0_0[31:31], simp432_0[0:0], simp432_0[1:1]);
  C3 I187 (simp441_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I188 (simp441_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I189 (simp441_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I190 (simp441_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  BUFF I191 (simp441_0[4:4], i_0r1[12:12]);
  C3 I192 (simp442_0[0:0], simp441_0[0:0], simp441_0[1:1], simp441_0[2:2]);
  C2 I193 (simp442_0[1:1], simp441_0[3:3], simp441_0[4:4]);
  C2 I194 (match0_0[32:32], simp442_0[0:0], simp442_0[1:1]);
  C3 I195 (simp451_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I196 (simp451_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I197 (simp451_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I198 (simp451_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  BUFF I199 (simp451_0[4:4], i_0r1[12:12]);
  C3 I200 (simp452_0[0:0], simp451_0[0:0], simp451_0[1:1], simp451_0[2:2]);
  C2 I201 (simp452_0[1:1], simp451_0[3:3], simp451_0[4:4]);
  C2 I202 (match0_0[33:33], simp452_0[0:0], simp452_0[1:1]);
  C3 I203 (simp461_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I204 (simp461_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I205 (simp461_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I206 (simp461_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C2 I207 (simp461_0[4:4], i_0r0[12:12], i_0r1[13:13]);
  C3 I208 (simp462_0[0:0], simp461_0[0:0], simp461_0[1:1], simp461_0[2:2]);
  C2 I209 (simp462_0[1:1], simp461_0[3:3], simp461_0[4:4]);
  C2 I210 (match0_0[34:34], simp462_0[0:0], simp462_0[1:1]);
  C3 I211 (simp471_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I212 (simp471_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I213 (simp471_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I214 (simp471_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C2 I215 (simp471_0[4:4], i_0r0[12:12], i_0r1[13:13]);
  C3 I216 (simp472_0[0:0], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  C2 I217 (simp472_0[1:1], simp471_0[3:3], simp471_0[4:4]);
  C2 I218 (match0_0[35:35], simp472_0[0:0], simp472_0[1:1]);
  C3 I219 (simp481_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I220 (simp481_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I221 (simp481_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I222 (simp481_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C2 I223 (simp481_0[4:4], i_0r0[12:12], i_0r1[13:13]);
  C3 I224 (simp482_0[0:0], simp481_0[0:0], simp481_0[1:1], simp481_0[2:2]);
  C2 I225 (simp482_0[1:1], simp481_0[3:3], simp481_0[4:4]);
  C2 I226 (match0_0[36:36], simp482_0[0:0], simp482_0[1:1]);
  C3 I227 (simp491_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I228 (simp491_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I229 (simp491_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I230 (simp491_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I231 (simp491_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r1[14:14]);
  C3 I232 (simp492_0[0:0], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  C2 I233 (simp492_0[1:1], simp491_0[3:3], simp491_0[4:4]);
  C2 I234 (match0_0[37:37], simp492_0[0:0], simp492_0[1:1]);
  C3 I235 (simp501_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I236 (simp501_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I237 (simp501_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I238 (simp501_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I239 (simp501_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r1[14:14]);
  C3 I240 (simp502_0[0:0], simp501_0[0:0], simp501_0[1:1], simp501_0[2:2]);
  C2 I241 (simp502_0[1:1], simp501_0[3:3], simp501_0[4:4]);
  C2 I242 (match0_0[38:38], simp502_0[0:0], simp502_0[1:1]);
  C3 I243 (simp511_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I244 (simp511_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I245 (simp511_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I246 (simp511_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I247 (simp511_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r1[14:14]);
  C3 I248 (simp512_0[0:0], simp511_0[0:0], simp511_0[1:1], simp511_0[2:2]);
  C2 I249 (simp512_0[1:1], simp511_0[3:3], simp511_0[4:4]);
  C2 I250 (match0_0[39:39], simp512_0[0:0], simp512_0[1:1]);
  C3 I251 (simp521_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I252 (simp521_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I253 (simp521_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I254 (simp521_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I255 (simp521_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  BUFF I256 (simp521_0[5:5], i_0r1[15:15]);
  C3 I257 (simp522_0[0:0], simp521_0[0:0], simp521_0[1:1], simp521_0[2:2]);
  C3 I258 (simp522_0[1:1], simp521_0[3:3], simp521_0[4:4], simp521_0[5:5]);
  C2 I259 (match0_0[40:40], simp522_0[0:0], simp522_0[1:1]);
  C3 I260 (simp531_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I261 (simp531_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I262 (simp531_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I263 (simp531_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I264 (simp531_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  BUFF I265 (simp531_0[5:5], i_0r1[15:15]);
  C3 I266 (simp532_0[0:0], simp531_0[0:0], simp531_0[1:1], simp531_0[2:2]);
  C3 I267 (simp532_0[1:1], simp531_0[3:3], simp531_0[4:4], simp531_0[5:5]);
  C2 I268 (match0_0[41:41], simp532_0[0:0], simp532_0[1:1]);
  C3 I269 (simp541_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I270 (simp541_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I271 (simp541_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I272 (simp541_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I273 (simp541_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  BUFF I274 (simp541_0[5:5], i_0r1[15:15]);
  C3 I275 (simp542_0[0:0], simp541_0[0:0], simp541_0[1:1], simp541_0[2:2]);
  C3 I276 (simp542_0[1:1], simp541_0[3:3], simp541_0[4:4], simp541_0[5:5]);
  C2 I277 (match0_0[42:42], simp542_0[0:0], simp542_0[1:1]);
  C3 I278 (simp551_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I279 (simp551_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I280 (simp551_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I281 (simp551_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I282 (simp551_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C2 I283 (simp551_0[5:5], i_0r0[15:15], i_0r1[16:16]);
  C3 I284 (simp552_0[0:0], simp551_0[0:0], simp551_0[1:1], simp551_0[2:2]);
  C3 I285 (simp552_0[1:1], simp551_0[3:3], simp551_0[4:4], simp551_0[5:5]);
  C2 I286 (match0_0[43:43], simp552_0[0:0], simp552_0[1:1]);
  C3 I287 (simp561_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I288 (simp561_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I289 (simp561_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I290 (simp561_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I291 (simp561_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C2 I292 (simp561_0[5:5], i_0r0[15:15], i_0r1[16:16]);
  C3 I293 (simp562_0[0:0], simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  C3 I294 (simp562_0[1:1], simp561_0[3:3], simp561_0[4:4], simp561_0[5:5]);
  C2 I295 (match0_0[44:44], simp562_0[0:0], simp562_0[1:1]);
  C3 I296 (simp571_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I297 (simp571_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I298 (simp571_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I299 (simp571_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I300 (simp571_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C2 I301 (simp571_0[5:5], i_0r0[15:15], i_0r1[16:16]);
  C3 I302 (simp572_0[0:0], simp571_0[0:0], simp571_0[1:1], simp571_0[2:2]);
  C3 I303 (simp572_0[1:1], simp571_0[3:3], simp571_0[4:4], simp571_0[5:5]);
  C2 I304 (match0_0[45:45], simp572_0[0:0], simp572_0[1:1]);
  C3 I305 (simp581_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I306 (simp581_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I307 (simp581_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I308 (simp581_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I309 (simp581_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I310 (simp581_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r1[17:17]);
  C3 I311 (simp582_0[0:0], simp581_0[0:0], simp581_0[1:1], simp581_0[2:2]);
  C3 I312 (simp582_0[1:1], simp581_0[3:3], simp581_0[4:4], simp581_0[5:5]);
  C2 I313 (match0_0[46:46], simp582_0[0:0], simp582_0[1:1]);
  C3 I314 (simp591_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I315 (simp591_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I316 (simp591_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I317 (simp591_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I318 (simp591_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I319 (simp591_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r1[17:17]);
  C3 I320 (simp592_0[0:0], simp591_0[0:0], simp591_0[1:1], simp591_0[2:2]);
  C3 I321 (simp592_0[1:1], simp591_0[3:3], simp591_0[4:4], simp591_0[5:5]);
  C2 I322 (match0_0[47:47], simp592_0[0:0], simp592_0[1:1]);
  C3 I323 (simp601_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I324 (simp601_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I325 (simp601_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I326 (simp601_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I327 (simp601_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I328 (simp601_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r1[17:17]);
  C3 I329 (simp602_0[0:0], simp601_0[0:0], simp601_0[1:1], simp601_0[2:2]);
  C3 I330 (simp602_0[1:1], simp601_0[3:3], simp601_0[4:4], simp601_0[5:5]);
  C2 I331 (match0_0[48:48], simp602_0[0:0], simp602_0[1:1]);
  C3 I332 (simp611_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I333 (simp611_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I334 (simp611_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I335 (simp611_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I336 (simp611_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I337 (simp611_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  BUFF I338 (simp611_0[6:6], i_0r1[18:18]);
  C3 I339 (simp612_0[0:0], simp611_0[0:0], simp611_0[1:1], simp611_0[2:2]);
  C3 I340 (simp612_0[1:1], simp611_0[3:3], simp611_0[4:4], simp611_0[5:5]);
  BUFF I341 (simp612_0[2:2], simp611_0[6:6]);
  C3 I342 (match0_0[49:49], simp612_0[0:0], simp612_0[1:1], simp612_0[2:2]);
  C3 I343 (simp621_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I344 (simp621_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I345 (simp621_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I346 (simp621_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I347 (simp621_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I348 (simp621_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  BUFF I349 (simp621_0[6:6], i_0r1[18:18]);
  C3 I350 (simp622_0[0:0], simp621_0[0:0], simp621_0[1:1], simp621_0[2:2]);
  C3 I351 (simp622_0[1:1], simp621_0[3:3], simp621_0[4:4], simp621_0[5:5]);
  BUFF I352 (simp622_0[2:2], simp621_0[6:6]);
  C3 I353 (match0_0[50:50], simp622_0[0:0], simp622_0[1:1], simp622_0[2:2]);
  C3 I354 (simp631_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I355 (simp631_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I356 (simp631_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I357 (simp631_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I358 (simp631_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I359 (simp631_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  BUFF I360 (simp631_0[6:6], i_0r1[18:18]);
  C3 I361 (simp632_0[0:0], simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  C3 I362 (simp632_0[1:1], simp631_0[3:3], simp631_0[4:4], simp631_0[5:5]);
  BUFF I363 (simp632_0[2:2], simp631_0[6:6]);
  C3 I364 (match0_0[51:51], simp632_0[0:0], simp632_0[1:1], simp632_0[2:2]);
  C3 I365 (simp641_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I366 (simp641_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I367 (simp641_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I368 (simp641_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I369 (simp641_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I370 (simp641_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C2 I371 (simp641_0[6:6], i_0r0[18:18], i_0r1[19:19]);
  C3 I372 (simp642_0[0:0], simp641_0[0:0], simp641_0[1:1], simp641_0[2:2]);
  C3 I373 (simp642_0[1:1], simp641_0[3:3], simp641_0[4:4], simp641_0[5:5]);
  BUFF I374 (simp642_0[2:2], simp641_0[6:6]);
  C3 I375 (match0_0[52:52], simp642_0[0:0], simp642_0[1:1], simp642_0[2:2]);
  C3 I376 (simp651_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I377 (simp651_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I378 (simp651_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I379 (simp651_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I380 (simp651_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I381 (simp651_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C2 I382 (simp651_0[6:6], i_0r0[18:18], i_0r1[19:19]);
  C3 I383 (simp652_0[0:0], simp651_0[0:0], simp651_0[1:1], simp651_0[2:2]);
  C3 I384 (simp652_0[1:1], simp651_0[3:3], simp651_0[4:4], simp651_0[5:5]);
  BUFF I385 (simp652_0[2:2], simp651_0[6:6]);
  C3 I386 (match0_0[53:53], simp652_0[0:0], simp652_0[1:1], simp652_0[2:2]);
  C3 I387 (simp661_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I388 (simp661_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I389 (simp661_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I390 (simp661_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I391 (simp661_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I392 (simp661_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C2 I393 (simp661_0[6:6], i_0r0[18:18], i_0r1[19:19]);
  C3 I394 (simp662_0[0:0], simp661_0[0:0], simp661_0[1:1], simp661_0[2:2]);
  C3 I395 (simp662_0[1:1], simp661_0[3:3], simp661_0[4:4], simp661_0[5:5]);
  BUFF I396 (simp662_0[2:2], simp661_0[6:6]);
  C3 I397 (match0_0[54:54], simp662_0[0:0], simp662_0[1:1], simp662_0[2:2]);
  C3 I398 (simp671_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I399 (simp671_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I400 (simp671_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I401 (simp671_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I402 (simp671_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I403 (simp671_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I404 (simp671_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r1[20:20]);
  C3 I405 (simp672_0[0:0], simp671_0[0:0], simp671_0[1:1], simp671_0[2:2]);
  C3 I406 (simp672_0[1:1], simp671_0[3:3], simp671_0[4:4], simp671_0[5:5]);
  BUFF I407 (simp672_0[2:2], simp671_0[6:6]);
  C3 I408 (match0_0[55:55], simp672_0[0:0], simp672_0[1:1], simp672_0[2:2]);
  C3 I409 (simp681_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I410 (simp681_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I411 (simp681_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I412 (simp681_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I413 (simp681_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I414 (simp681_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I415 (simp681_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r1[20:20]);
  C3 I416 (simp682_0[0:0], simp681_0[0:0], simp681_0[1:1], simp681_0[2:2]);
  C3 I417 (simp682_0[1:1], simp681_0[3:3], simp681_0[4:4], simp681_0[5:5]);
  BUFF I418 (simp682_0[2:2], simp681_0[6:6]);
  C3 I419 (match0_0[56:56], simp682_0[0:0], simp682_0[1:1], simp682_0[2:2]);
  C3 I420 (simp691_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I421 (simp691_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I422 (simp691_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I423 (simp691_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I424 (simp691_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I425 (simp691_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I426 (simp691_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r1[20:20]);
  C3 I427 (simp692_0[0:0], simp691_0[0:0], simp691_0[1:1], simp691_0[2:2]);
  C3 I428 (simp692_0[1:1], simp691_0[3:3], simp691_0[4:4], simp691_0[5:5]);
  BUFF I429 (simp692_0[2:2], simp691_0[6:6]);
  C3 I430 (match0_0[57:57], simp692_0[0:0], simp692_0[1:1], simp692_0[2:2]);
  C3 I431 (simp701_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I432 (simp701_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I433 (simp701_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I434 (simp701_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I435 (simp701_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I436 (simp701_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I437 (simp701_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  BUFF I438 (simp701_0[7:7], i_0r1[21:21]);
  C3 I439 (simp702_0[0:0], simp701_0[0:0], simp701_0[1:1], simp701_0[2:2]);
  C3 I440 (simp702_0[1:1], simp701_0[3:3], simp701_0[4:4], simp701_0[5:5]);
  C2 I441 (simp702_0[2:2], simp701_0[6:6], simp701_0[7:7]);
  C3 I442 (match0_0[58:58], simp702_0[0:0], simp702_0[1:1], simp702_0[2:2]);
  C3 I443 (simp711_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I444 (simp711_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I445 (simp711_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I446 (simp711_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I447 (simp711_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I448 (simp711_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I449 (simp711_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  BUFF I450 (simp711_0[7:7], i_0r1[21:21]);
  C3 I451 (simp712_0[0:0], simp711_0[0:0], simp711_0[1:1], simp711_0[2:2]);
  C3 I452 (simp712_0[1:1], simp711_0[3:3], simp711_0[4:4], simp711_0[5:5]);
  C2 I453 (simp712_0[2:2], simp711_0[6:6], simp711_0[7:7]);
  C3 I454 (match0_0[59:59], simp712_0[0:0], simp712_0[1:1], simp712_0[2:2]);
  C3 I455 (simp721_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I456 (simp721_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I457 (simp721_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I458 (simp721_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I459 (simp721_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I460 (simp721_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I461 (simp721_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  BUFF I462 (simp721_0[7:7], i_0r1[21:21]);
  C3 I463 (simp722_0[0:0], simp721_0[0:0], simp721_0[1:1], simp721_0[2:2]);
  C3 I464 (simp722_0[1:1], simp721_0[3:3], simp721_0[4:4], simp721_0[5:5]);
  C2 I465 (simp722_0[2:2], simp721_0[6:6], simp721_0[7:7]);
  C3 I466 (match0_0[60:60], simp722_0[0:0], simp722_0[1:1], simp722_0[2:2]);
  C3 I467 (simp731_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I468 (simp731_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I469 (simp731_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I470 (simp731_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I471 (simp731_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I472 (simp731_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I473 (simp731_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C2 I474 (simp731_0[7:7], i_0r0[21:21], i_0r1[22:22]);
  C3 I475 (simp732_0[0:0], simp731_0[0:0], simp731_0[1:1], simp731_0[2:2]);
  C3 I476 (simp732_0[1:1], simp731_0[3:3], simp731_0[4:4], simp731_0[5:5]);
  C2 I477 (simp732_0[2:2], simp731_0[6:6], simp731_0[7:7]);
  C3 I478 (match0_0[61:61], simp732_0[0:0], simp732_0[1:1], simp732_0[2:2]);
  C3 I479 (simp741_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I480 (simp741_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I481 (simp741_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I482 (simp741_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I483 (simp741_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I484 (simp741_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I485 (simp741_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C2 I486 (simp741_0[7:7], i_0r0[21:21], i_0r1[22:22]);
  C3 I487 (simp742_0[0:0], simp741_0[0:0], simp741_0[1:1], simp741_0[2:2]);
  C3 I488 (simp742_0[1:1], simp741_0[3:3], simp741_0[4:4], simp741_0[5:5]);
  C2 I489 (simp742_0[2:2], simp741_0[6:6], simp741_0[7:7]);
  C3 I490 (match0_0[62:62], simp742_0[0:0], simp742_0[1:1], simp742_0[2:2]);
  C3 I491 (simp751_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I492 (simp751_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I493 (simp751_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I494 (simp751_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I495 (simp751_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I496 (simp751_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I497 (simp751_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C2 I498 (simp751_0[7:7], i_0r0[21:21], i_0r1[22:22]);
  C3 I499 (simp752_0[0:0], simp751_0[0:0], simp751_0[1:1], simp751_0[2:2]);
  C3 I500 (simp752_0[1:1], simp751_0[3:3], simp751_0[4:4], simp751_0[5:5]);
  C2 I501 (simp752_0[2:2], simp751_0[6:6], simp751_0[7:7]);
  C3 I502 (match0_0[63:63], simp752_0[0:0], simp752_0[1:1], simp752_0[2:2]);
  C3 I503 (simp761_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I504 (simp761_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I505 (simp761_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I506 (simp761_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I507 (simp761_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I508 (simp761_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I509 (simp761_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I510 (simp761_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r1[23:23]);
  C3 I511 (simp762_0[0:0], simp761_0[0:0], simp761_0[1:1], simp761_0[2:2]);
  C3 I512 (simp762_0[1:1], simp761_0[3:3], simp761_0[4:4], simp761_0[5:5]);
  C2 I513 (simp762_0[2:2], simp761_0[6:6], simp761_0[7:7]);
  C3 I514 (match0_0[64:64], simp762_0[0:0], simp762_0[1:1], simp762_0[2:2]);
  C3 I515 (simp771_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I516 (simp771_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I517 (simp771_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I518 (simp771_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I519 (simp771_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I520 (simp771_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I521 (simp771_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I522 (simp771_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r1[23:23]);
  C3 I523 (simp772_0[0:0], simp771_0[0:0], simp771_0[1:1], simp771_0[2:2]);
  C3 I524 (simp772_0[1:1], simp771_0[3:3], simp771_0[4:4], simp771_0[5:5]);
  C2 I525 (simp772_0[2:2], simp771_0[6:6], simp771_0[7:7]);
  C3 I526 (match0_0[65:65], simp772_0[0:0], simp772_0[1:1], simp772_0[2:2]);
  C3 I527 (simp781_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I528 (simp781_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I529 (simp781_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I530 (simp781_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I531 (simp781_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I532 (simp781_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I533 (simp781_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I534 (simp781_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r1[23:23]);
  C3 I535 (simp782_0[0:0], simp781_0[0:0], simp781_0[1:1], simp781_0[2:2]);
  C3 I536 (simp782_0[1:1], simp781_0[3:3], simp781_0[4:4], simp781_0[5:5]);
  C2 I537 (simp782_0[2:2], simp781_0[6:6], simp781_0[7:7]);
  C3 I538 (match0_0[66:66], simp782_0[0:0], simp782_0[1:1], simp782_0[2:2]);
  C3 I539 (simp791_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I540 (simp791_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I541 (simp791_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I542 (simp791_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I543 (simp791_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I544 (simp791_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I545 (simp791_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I546 (simp791_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  BUFF I547 (simp791_0[8:8], i_0r1[24:24]);
  C3 I548 (simp792_0[0:0], simp791_0[0:0], simp791_0[1:1], simp791_0[2:2]);
  C3 I549 (simp792_0[1:1], simp791_0[3:3], simp791_0[4:4], simp791_0[5:5]);
  C3 I550 (simp792_0[2:2], simp791_0[6:6], simp791_0[7:7], simp791_0[8:8]);
  C3 I551 (match0_0[67:67], simp792_0[0:0], simp792_0[1:1], simp792_0[2:2]);
  C3 I552 (simp801_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I553 (simp801_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I554 (simp801_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I555 (simp801_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I556 (simp801_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I557 (simp801_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I558 (simp801_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I559 (simp801_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  BUFF I560 (simp801_0[8:8], i_0r1[24:24]);
  C3 I561 (simp802_0[0:0], simp801_0[0:0], simp801_0[1:1], simp801_0[2:2]);
  C3 I562 (simp802_0[1:1], simp801_0[3:3], simp801_0[4:4], simp801_0[5:5]);
  C3 I563 (simp802_0[2:2], simp801_0[6:6], simp801_0[7:7], simp801_0[8:8]);
  C3 I564 (match0_0[68:68], simp802_0[0:0], simp802_0[1:1], simp802_0[2:2]);
  C3 I565 (simp811_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I566 (simp811_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I567 (simp811_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I568 (simp811_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I569 (simp811_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I570 (simp811_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I571 (simp811_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I572 (simp811_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  BUFF I573 (simp811_0[8:8], i_0r1[24:24]);
  C3 I574 (simp812_0[0:0], simp811_0[0:0], simp811_0[1:1], simp811_0[2:2]);
  C3 I575 (simp812_0[1:1], simp811_0[3:3], simp811_0[4:4], simp811_0[5:5]);
  C3 I576 (simp812_0[2:2], simp811_0[6:6], simp811_0[7:7], simp811_0[8:8]);
  C3 I577 (match0_0[69:69], simp812_0[0:0], simp812_0[1:1], simp812_0[2:2]);
  C3 I578 (simp821_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I579 (simp821_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I580 (simp821_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I581 (simp821_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I582 (simp821_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I583 (simp821_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I584 (simp821_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I585 (simp821_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C2 I586 (simp821_0[8:8], i_0r0[24:24], i_0r1[25:25]);
  C3 I587 (simp822_0[0:0], simp821_0[0:0], simp821_0[1:1], simp821_0[2:2]);
  C3 I588 (simp822_0[1:1], simp821_0[3:3], simp821_0[4:4], simp821_0[5:5]);
  C3 I589 (simp822_0[2:2], simp821_0[6:6], simp821_0[7:7], simp821_0[8:8]);
  C3 I590 (match0_0[70:70], simp822_0[0:0], simp822_0[1:1], simp822_0[2:2]);
  C3 I591 (simp831_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I592 (simp831_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I593 (simp831_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I594 (simp831_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I595 (simp831_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I596 (simp831_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I597 (simp831_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I598 (simp831_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C2 I599 (simp831_0[8:8], i_0r0[24:24], i_0r1[25:25]);
  C3 I600 (simp832_0[0:0], simp831_0[0:0], simp831_0[1:1], simp831_0[2:2]);
  C3 I601 (simp832_0[1:1], simp831_0[3:3], simp831_0[4:4], simp831_0[5:5]);
  C3 I602 (simp832_0[2:2], simp831_0[6:6], simp831_0[7:7], simp831_0[8:8]);
  C3 I603 (match0_0[71:71], simp832_0[0:0], simp832_0[1:1], simp832_0[2:2]);
  C3 I604 (simp841_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I605 (simp841_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I606 (simp841_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I607 (simp841_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I608 (simp841_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I609 (simp841_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I610 (simp841_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I611 (simp841_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C2 I612 (simp841_0[8:8], i_0r0[24:24], i_0r1[25:25]);
  C3 I613 (simp842_0[0:0], simp841_0[0:0], simp841_0[1:1], simp841_0[2:2]);
  C3 I614 (simp842_0[1:1], simp841_0[3:3], simp841_0[4:4], simp841_0[5:5]);
  C3 I615 (simp842_0[2:2], simp841_0[6:6], simp841_0[7:7], simp841_0[8:8]);
  C3 I616 (match0_0[72:72], simp842_0[0:0], simp842_0[1:1], simp842_0[2:2]);
  C3 I617 (simp851_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I618 (simp851_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I619 (simp851_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I620 (simp851_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I621 (simp851_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I622 (simp851_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I623 (simp851_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I624 (simp851_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I625 (simp851_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r1[26:26]);
  C3 I626 (simp852_0[0:0], simp851_0[0:0], simp851_0[1:1], simp851_0[2:2]);
  C3 I627 (simp852_0[1:1], simp851_0[3:3], simp851_0[4:4], simp851_0[5:5]);
  C3 I628 (simp852_0[2:2], simp851_0[6:6], simp851_0[7:7], simp851_0[8:8]);
  C3 I629 (match0_0[73:73], simp852_0[0:0], simp852_0[1:1], simp852_0[2:2]);
  C3 I630 (simp861_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I631 (simp861_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I632 (simp861_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I633 (simp861_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I634 (simp861_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I635 (simp861_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I636 (simp861_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I637 (simp861_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I638 (simp861_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r1[26:26]);
  C3 I639 (simp862_0[0:0], simp861_0[0:0], simp861_0[1:1], simp861_0[2:2]);
  C3 I640 (simp862_0[1:1], simp861_0[3:3], simp861_0[4:4], simp861_0[5:5]);
  C3 I641 (simp862_0[2:2], simp861_0[6:6], simp861_0[7:7], simp861_0[8:8]);
  C3 I642 (match0_0[74:74], simp862_0[0:0], simp862_0[1:1], simp862_0[2:2]);
  C3 I643 (simp871_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I644 (simp871_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I645 (simp871_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I646 (simp871_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I647 (simp871_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I648 (simp871_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I649 (simp871_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I650 (simp871_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I651 (simp871_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r1[26:26]);
  C3 I652 (simp872_0[0:0], simp871_0[0:0], simp871_0[1:1], simp871_0[2:2]);
  C3 I653 (simp872_0[1:1], simp871_0[3:3], simp871_0[4:4], simp871_0[5:5]);
  C3 I654 (simp872_0[2:2], simp871_0[6:6], simp871_0[7:7], simp871_0[8:8]);
  C3 I655 (match0_0[75:75], simp872_0[0:0], simp872_0[1:1], simp872_0[2:2]);
  C3 I656 (simp881_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I657 (simp881_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I658 (simp881_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I659 (simp881_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I660 (simp881_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I661 (simp881_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I662 (simp881_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I663 (simp881_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I664 (simp881_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  BUFF I665 (simp881_0[9:9], i_0r1[27:27]);
  C3 I666 (simp882_0[0:0], simp881_0[0:0], simp881_0[1:1], simp881_0[2:2]);
  C3 I667 (simp882_0[1:1], simp881_0[3:3], simp881_0[4:4], simp881_0[5:5]);
  C3 I668 (simp882_0[2:2], simp881_0[6:6], simp881_0[7:7], simp881_0[8:8]);
  BUFF I669 (simp882_0[3:3], simp881_0[9:9]);
  C3 I670 (simp883_0[0:0], simp882_0[0:0], simp882_0[1:1], simp882_0[2:2]);
  BUFF I671 (simp883_0[1:1], simp882_0[3:3]);
  C2 I672 (match0_0[76:76], simp883_0[0:0], simp883_0[1:1]);
  C3 I673 (simp891_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I674 (simp891_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I675 (simp891_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I676 (simp891_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I677 (simp891_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I678 (simp891_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I679 (simp891_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I680 (simp891_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I681 (simp891_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  BUFF I682 (simp891_0[9:9], i_0r1[27:27]);
  C3 I683 (simp892_0[0:0], simp891_0[0:0], simp891_0[1:1], simp891_0[2:2]);
  C3 I684 (simp892_0[1:1], simp891_0[3:3], simp891_0[4:4], simp891_0[5:5]);
  C3 I685 (simp892_0[2:2], simp891_0[6:6], simp891_0[7:7], simp891_0[8:8]);
  BUFF I686 (simp892_0[3:3], simp891_0[9:9]);
  C3 I687 (simp893_0[0:0], simp892_0[0:0], simp892_0[1:1], simp892_0[2:2]);
  BUFF I688 (simp893_0[1:1], simp892_0[3:3]);
  C2 I689 (match0_0[77:77], simp893_0[0:0], simp893_0[1:1]);
  C3 I690 (simp901_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I691 (simp901_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I692 (simp901_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I693 (simp901_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I694 (simp901_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I695 (simp901_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I696 (simp901_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I697 (simp901_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I698 (simp901_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  BUFF I699 (simp901_0[9:9], i_0r1[27:27]);
  C3 I700 (simp902_0[0:0], simp901_0[0:0], simp901_0[1:1], simp901_0[2:2]);
  C3 I701 (simp902_0[1:1], simp901_0[3:3], simp901_0[4:4], simp901_0[5:5]);
  C3 I702 (simp902_0[2:2], simp901_0[6:6], simp901_0[7:7], simp901_0[8:8]);
  BUFF I703 (simp902_0[3:3], simp901_0[9:9]);
  C3 I704 (simp903_0[0:0], simp902_0[0:0], simp902_0[1:1], simp902_0[2:2]);
  BUFF I705 (simp903_0[1:1], simp902_0[3:3]);
  C2 I706 (match0_0[78:78], simp903_0[0:0], simp903_0[1:1]);
  C3 I707 (simp911_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I708 (simp911_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I709 (simp911_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I710 (simp911_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I711 (simp911_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I712 (simp911_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I713 (simp911_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I714 (simp911_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I715 (simp911_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C2 I716 (simp911_0[9:9], i_0r0[27:27], i_0r1[28:28]);
  C3 I717 (simp912_0[0:0], simp911_0[0:0], simp911_0[1:1], simp911_0[2:2]);
  C3 I718 (simp912_0[1:1], simp911_0[3:3], simp911_0[4:4], simp911_0[5:5]);
  C3 I719 (simp912_0[2:2], simp911_0[6:6], simp911_0[7:7], simp911_0[8:8]);
  BUFF I720 (simp912_0[3:3], simp911_0[9:9]);
  C3 I721 (simp913_0[0:0], simp912_0[0:0], simp912_0[1:1], simp912_0[2:2]);
  BUFF I722 (simp913_0[1:1], simp912_0[3:3]);
  C2 I723 (match0_0[79:79], simp913_0[0:0], simp913_0[1:1]);
  C3 I724 (simp921_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I725 (simp921_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I726 (simp921_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I727 (simp921_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I728 (simp921_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I729 (simp921_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I730 (simp921_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I731 (simp921_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I732 (simp921_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C2 I733 (simp921_0[9:9], i_0r0[27:27], i_0r1[28:28]);
  C3 I734 (simp922_0[0:0], simp921_0[0:0], simp921_0[1:1], simp921_0[2:2]);
  C3 I735 (simp922_0[1:1], simp921_0[3:3], simp921_0[4:4], simp921_0[5:5]);
  C3 I736 (simp922_0[2:2], simp921_0[6:6], simp921_0[7:7], simp921_0[8:8]);
  BUFF I737 (simp922_0[3:3], simp921_0[9:9]);
  C3 I738 (simp923_0[0:0], simp922_0[0:0], simp922_0[1:1], simp922_0[2:2]);
  BUFF I739 (simp923_0[1:1], simp922_0[3:3]);
  C2 I740 (match0_0[80:80], simp923_0[0:0], simp923_0[1:1]);
  C3 I741 (simp931_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I742 (simp931_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I743 (simp931_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I744 (simp931_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I745 (simp931_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I746 (simp931_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I747 (simp931_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I748 (simp931_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I749 (simp931_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C2 I750 (simp931_0[9:9], i_0r0[27:27], i_0r1[28:28]);
  C3 I751 (simp932_0[0:0], simp931_0[0:0], simp931_0[1:1], simp931_0[2:2]);
  C3 I752 (simp932_0[1:1], simp931_0[3:3], simp931_0[4:4], simp931_0[5:5]);
  C3 I753 (simp932_0[2:2], simp931_0[6:6], simp931_0[7:7], simp931_0[8:8]);
  BUFF I754 (simp932_0[3:3], simp931_0[9:9]);
  C3 I755 (simp933_0[0:0], simp932_0[0:0], simp932_0[1:1], simp932_0[2:2]);
  BUFF I756 (simp933_0[1:1], simp932_0[3:3]);
  C2 I757 (match0_0[81:81], simp933_0[0:0], simp933_0[1:1]);
  C3 I758 (simp941_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I759 (simp941_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I760 (simp941_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I761 (simp941_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I762 (simp941_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I763 (simp941_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I764 (simp941_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I765 (simp941_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I766 (simp941_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I767 (simp941_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r1[29:29]);
  C3 I768 (simp942_0[0:0], simp941_0[0:0], simp941_0[1:1], simp941_0[2:2]);
  C3 I769 (simp942_0[1:1], simp941_0[3:3], simp941_0[4:4], simp941_0[5:5]);
  C3 I770 (simp942_0[2:2], simp941_0[6:6], simp941_0[7:7], simp941_0[8:8]);
  BUFF I771 (simp942_0[3:3], simp941_0[9:9]);
  C3 I772 (simp943_0[0:0], simp942_0[0:0], simp942_0[1:1], simp942_0[2:2]);
  BUFF I773 (simp943_0[1:1], simp942_0[3:3]);
  C2 I774 (match0_0[82:82], simp943_0[0:0], simp943_0[1:1]);
  C3 I775 (simp951_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I776 (simp951_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I777 (simp951_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I778 (simp951_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I779 (simp951_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I780 (simp951_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I781 (simp951_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I782 (simp951_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I783 (simp951_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I784 (simp951_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r1[29:29]);
  C3 I785 (simp952_0[0:0], simp951_0[0:0], simp951_0[1:1], simp951_0[2:2]);
  C3 I786 (simp952_0[1:1], simp951_0[3:3], simp951_0[4:4], simp951_0[5:5]);
  C3 I787 (simp952_0[2:2], simp951_0[6:6], simp951_0[7:7], simp951_0[8:8]);
  BUFF I788 (simp952_0[3:3], simp951_0[9:9]);
  C3 I789 (simp953_0[0:0], simp952_0[0:0], simp952_0[1:1], simp952_0[2:2]);
  BUFF I790 (simp953_0[1:1], simp952_0[3:3]);
  C2 I791 (match0_0[83:83], simp953_0[0:0], simp953_0[1:1]);
  C3 I792 (simp961_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I793 (simp961_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I794 (simp961_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I795 (simp961_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I796 (simp961_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I797 (simp961_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I798 (simp961_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I799 (simp961_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I800 (simp961_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I801 (simp961_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r1[29:29]);
  C3 I802 (simp962_0[0:0], simp961_0[0:0], simp961_0[1:1], simp961_0[2:2]);
  C3 I803 (simp962_0[1:1], simp961_0[3:3], simp961_0[4:4], simp961_0[5:5]);
  C3 I804 (simp962_0[2:2], simp961_0[6:6], simp961_0[7:7], simp961_0[8:8]);
  BUFF I805 (simp962_0[3:3], simp961_0[9:9]);
  C3 I806 (simp963_0[0:0], simp962_0[0:0], simp962_0[1:1], simp962_0[2:2]);
  BUFF I807 (simp963_0[1:1], simp962_0[3:3]);
  C2 I808 (match0_0[84:84], simp963_0[0:0], simp963_0[1:1]);
  C3 I809 (simp971_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I810 (simp971_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I811 (simp971_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I812 (simp971_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I813 (simp971_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I814 (simp971_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I815 (simp971_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I816 (simp971_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I817 (simp971_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I818 (simp971_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  BUFF I819 (simp971_0[10:10], i_0r1[30:30]);
  C3 I820 (simp972_0[0:0], simp971_0[0:0], simp971_0[1:1], simp971_0[2:2]);
  C3 I821 (simp972_0[1:1], simp971_0[3:3], simp971_0[4:4], simp971_0[5:5]);
  C3 I822 (simp972_0[2:2], simp971_0[6:6], simp971_0[7:7], simp971_0[8:8]);
  C2 I823 (simp972_0[3:3], simp971_0[9:9], simp971_0[10:10]);
  C3 I824 (simp973_0[0:0], simp972_0[0:0], simp972_0[1:1], simp972_0[2:2]);
  BUFF I825 (simp973_0[1:1], simp972_0[3:3]);
  C2 I826 (match0_0[85:85], simp973_0[0:0], simp973_0[1:1]);
  C3 I827 (simp981_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I828 (simp981_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I829 (simp981_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I830 (simp981_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I831 (simp981_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I832 (simp981_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I833 (simp981_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I834 (simp981_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I835 (simp981_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I836 (simp981_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  BUFF I837 (simp981_0[10:10], i_0r1[30:30]);
  C3 I838 (simp982_0[0:0], simp981_0[0:0], simp981_0[1:1], simp981_0[2:2]);
  C3 I839 (simp982_0[1:1], simp981_0[3:3], simp981_0[4:4], simp981_0[5:5]);
  C3 I840 (simp982_0[2:2], simp981_0[6:6], simp981_0[7:7], simp981_0[8:8]);
  C2 I841 (simp982_0[3:3], simp981_0[9:9], simp981_0[10:10]);
  C3 I842 (simp983_0[0:0], simp982_0[0:0], simp982_0[1:1], simp982_0[2:2]);
  BUFF I843 (simp983_0[1:1], simp982_0[3:3]);
  C2 I844 (match0_0[86:86], simp983_0[0:0], simp983_0[1:1]);
  C3 I845 (simp991_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I846 (simp991_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I847 (simp991_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I848 (simp991_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I849 (simp991_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I850 (simp991_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I851 (simp991_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I852 (simp991_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I853 (simp991_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I854 (simp991_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  BUFF I855 (simp991_0[10:10], i_0r1[30:30]);
  C3 I856 (simp992_0[0:0], simp991_0[0:0], simp991_0[1:1], simp991_0[2:2]);
  C3 I857 (simp992_0[1:1], simp991_0[3:3], simp991_0[4:4], simp991_0[5:5]);
  C3 I858 (simp992_0[2:2], simp991_0[6:6], simp991_0[7:7], simp991_0[8:8]);
  C2 I859 (simp992_0[3:3], simp991_0[9:9], simp991_0[10:10]);
  C3 I860 (simp993_0[0:0], simp992_0[0:0], simp992_0[1:1], simp992_0[2:2]);
  BUFF I861 (simp993_0[1:1], simp992_0[3:3]);
  C2 I862 (match0_0[87:87], simp993_0[0:0], simp993_0[1:1]);
  C3 I863 (simp1001_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I864 (simp1001_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I865 (simp1001_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I866 (simp1001_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I867 (simp1001_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I868 (simp1001_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I869 (simp1001_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I870 (simp1001_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I871 (simp1001_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I872 (simp1001_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  C2 I873 (simp1001_0[10:10], i_0r0[30:30], i_0r1[31:31]);
  C3 I874 (simp1002_0[0:0], simp1001_0[0:0], simp1001_0[1:1], simp1001_0[2:2]);
  C3 I875 (simp1002_0[1:1], simp1001_0[3:3], simp1001_0[4:4], simp1001_0[5:5]);
  C3 I876 (simp1002_0[2:2], simp1001_0[6:6], simp1001_0[7:7], simp1001_0[8:8]);
  C2 I877 (simp1002_0[3:3], simp1001_0[9:9], simp1001_0[10:10]);
  C3 I878 (simp1003_0[0:0], simp1002_0[0:0], simp1002_0[1:1], simp1002_0[2:2]);
  BUFF I879 (simp1003_0[1:1], simp1002_0[3:3]);
  C2 I880 (match0_0[88:88], simp1003_0[0:0], simp1003_0[1:1]);
  C3 I881 (simp1011_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I882 (simp1011_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I883 (simp1011_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I884 (simp1011_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I885 (simp1011_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I886 (simp1011_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I887 (simp1011_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I888 (simp1011_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I889 (simp1011_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I890 (simp1011_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  C2 I891 (simp1011_0[10:10], i_0r0[30:30], i_0r1[31:31]);
  C3 I892 (simp1012_0[0:0], simp1011_0[0:0], simp1011_0[1:1], simp1011_0[2:2]);
  C3 I893 (simp1012_0[1:1], simp1011_0[3:3], simp1011_0[4:4], simp1011_0[5:5]);
  C3 I894 (simp1012_0[2:2], simp1011_0[6:6], simp1011_0[7:7], simp1011_0[8:8]);
  C2 I895 (simp1012_0[3:3], simp1011_0[9:9], simp1011_0[10:10]);
  C3 I896 (simp1013_0[0:0], simp1012_0[0:0], simp1012_0[1:1], simp1012_0[2:2]);
  BUFF I897 (simp1013_0[1:1], simp1012_0[3:3]);
  C2 I898 (match0_0[89:89], simp1013_0[0:0], simp1013_0[1:1]);
  C3 I899 (simp1021_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I900 (simp1021_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I901 (simp1021_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I902 (simp1021_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I903 (simp1021_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I904 (simp1021_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I905 (simp1021_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I906 (simp1021_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I907 (simp1021_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I908 (simp1021_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  C2 I909 (simp1021_0[10:10], i_0r0[30:30], i_0r1[31:31]);
  C3 I910 (simp1022_0[0:0], simp1021_0[0:0], simp1021_0[1:1], simp1021_0[2:2]);
  C3 I911 (simp1022_0[1:1], simp1021_0[3:3], simp1021_0[4:4], simp1021_0[5:5]);
  C3 I912 (simp1022_0[2:2], simp1021_0[6:6], simp1021_0[7:7], simp1021_0[8:8]);
  C2 I913 (simp1022_0[3:3], simp1021_0[9:9], simp1021_0[10:10]);
  C3 I914 (simp1023_0[0:0], simp1022_0[0:0], simp1022_0[1:1], simp1022_0[2:2]);
  BUFF I915 (simp1023_0[1:1], simp1022_0[3:3]);
  C2 I916 (match0_0[90:90], simp1023_0[0:0], simp1023_0[1:1]);
  BUFF I917 (sel_1, match1_0);
  C3 I918 (simp1051_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I919 (simp1051_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I920 (simp1051_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I921 (simp1051_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I922 (simp1051_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I923 (simp1051_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I924 (simp1051_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I925 (simp1051_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I926 (simp1051_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I927 (simp1051_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  C2 I928 (simp1051_0[10:10], i_0r0[30:30], i_0r0[31:31]);
  C3 I929 (simp1052_0[0:0], simp1051_0[0:0], simp1051_0[1:1], simp1051_0[2:2]);
  C3 I930 (simp1052_0[1:1], simp1051_0[3:3], simp1051_0[4:4], simp1051_0[5:5]);
  C3 I931 (simp1052_0[2:2], simp1051_0[6:6], simp1051_0[7:7], simp1051_0[8:8]);
  C2 I932 (simp1052_0[3:3], simp1051_0[9:9], simp1051_0[10:10]);
  C3 I933 (simp1053_0[0:0], simp1052_0[0:0], simp1052_0[1:1], simp1052_0[2:2]);
  BUFF I934 (simp1053_0[1:1], simp1052_0[3:3]);
  C2 I935 (match1_0, simp1053_0[0:0], simp1053_0[1:1]);
  BUFF I936 (sel_2, match2_0);
  C3 I937 (simp1081_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I938 (simp1081_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I939 (simp1081_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I940 (simp1081_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I941 (simp1081_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I942 (simp1081_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I943 (simp1081_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I944 (simp1081_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I945 (simp1081_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I946 (simp1081_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  C2 I947 (simp1081_0[10:10], i_0r0[30:30], i_0r0[31:31]);
  C3 I948 (simp1082_0[0:0], simp1081_0[0:0], simp1081_0[1:1], simp1081_0[2:2]);
  C3 I949 (simp1082_0[1:1], simp1081_0[3:3], simp1081_0[4:4], simp1081_0[5:5]);
  C3 I950 (simp1082_0[2:2], simp1081_0[6:6], simp1081_0[7:7], simp1081_0[8:8]);
  C2 I951 (simp1082_0[3:3], simp1081_0[9:9], simp1081_0[10:10]);
  C3 I952 (simp1083_0[0:0], simp1082_0[0:0], simp1082_0[1:1], simp1082_0[2:2]);
  BUFF I953 (simp1083_0[1:1], simp1082_0[3:3]);
  C2 I954 (match2_0, simp1083_0[0:0], simp1083_0[1:1]);
  BUFF I955 (sel_3, match3_0);
  C3 I956 (simp1111_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I957 (simp1111_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I958 (simp1111_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C3 I959 (simp1111_0[3:3], i_0r0[9:9], i_0r0[10:10], i_0r0[11:11]);
  C3 I960 (simp1111_0[4:4], i_0r0[12:12], i_0r0[13:13], i_0r0[14:14]);
  C3 I961 (simp1111_0[5:5], i_0r0[15:15], i_0r0[16:16], i_0r0[17:17]);
  C3 I962 (simp1111_0[6:6], i_0r0[18:18], i_0r0[19:19], i_0r0[20:20]);
  C3 I963 (simp1111_0[7:7], i_0r0[21:21], i_0r0[22:22], i_0r0[23:23]);
  C3 I964 (simp1111_0[8:8], i_0r0[24:24], i_0r0[25:25], i_0r0[26:26]);
  C3 I965 (simp1111_0[9:9], i_0r0[27:27], i_0r0[28:28], i_0r0[29:29]);
  C2 I966 (simp1111_0[10:10], i_0r0[30:30], i_0r0[31:31]);
  C3 I967 (simp1112_0[0:0], simp1111_0[0:0], simp1111_0[1:1], simp1111_0[2:2]);
  C3 I968 (simp1112_0[1:1], simp1111_0[3:3], simp1111_0[4:4], simp1111_0[5:5]);
  C3 I969 (simp1112_0[2:2], simp1111_0[6:6], simp1111_0[7:7], simp1111_0[8:8]);
  C2 I970 (simp1112_0[3:3], simp1111_0[9:9], simp1111_0[10:10]);
  C3 I971 (simp1113_0[0:0], simp1112_0[0:0], simp1112_0[1:1], simp1112_0[2:2]);
  BUFF I972 (simp1113_0[1:1], simp1112_0[3:3]);
  C2 I973 (match3_0, simp1113_0[0:0], simp1113_0[1:1]);
  C2 I974 (gsel_0, sel_0, icomplete_0);
  C2 I975 (gsel_1, sel_1, icomplete_0);
  C2 I976 (gsel_2, sel_2, icomplete_0);
  C2 I977 (gsel_3, sel_3, icomplete_0);
  OR2 I978 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I979 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I980 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I981 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I982 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I983 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I984 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I985 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I986 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I987 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I988 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I989 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I990 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I991 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I992 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I993 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I994 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I995 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I996 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I997 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I998 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I999 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I1000 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I1001 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I1002 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I1003 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I1004 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I1005 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I1006 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I1007 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I1008 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I1009 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I1010 (simp1491_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I1011 (simp1491_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I1012 (simp1491_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I1013 (simp1491_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I1014 (simp1491_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I1015 (simp1491_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I1016 (simp1491_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I1017 (simp1491_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I1018 (simp1491_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I1019 (simp1491_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C2 I1020 (simp1491_0[10:10], comp_0[30:30], comp_0[31:31]);
  C3 I1021 (simp1492_0[0:0], simp1491_0[0:0], simp1491_0[1:1], simp1491_0[2:2]);
  C3 I1022 (simp1492_0[1:1], simp1491_0[3:3], simp1491_0[4:4], simp1491_0[5:5]);
  C3 I1023 (simp1492_0[2:2], simp1491_0[6:6], simp1491_0[7:7], simp1491_0[8:8]);
  C2 I1024 (simp1492_0[3:3], simp1491_0[9:9], simp1491_0[10:10]);
  C3 I1025 (simp1493_0[0:0], simp1492_0[0:0], simp1492_0[1:1], simp1492_0[2:2]);
  BUFF I1026 (simp1493_0[1:1], simp1492_0[3:3]);
  C2 I1027 (icomplete_0, simp1493_0[0:0], simp1493_0[1:1]);
  BUFF I1028 (o_0r, gsel_0);
  BUFF I1029 (o_1r, gsel_1);
  BUFF I1030 (o_2r, gsel_2);
  BUFF I1031 (o_3r, gsel_3);
  NOR3 I1032 (simp1541_0[0:0], o_0a, o_1a, o_2a);
  INV I1033 (simp1541_0[1:1], o_3a);
  NAND2 I1034 (oack_0, simp1541_0[0:0], simp1541_0[1:1]);
  C2 I1035 (i_0a, oack_0, icomplete_0);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0] [One 0,Many [0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  input reset;
  wire [1:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  C3 I5 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C2 I6 (simp11_0[1:1], o_3a, o_4a);
  C2 I7 (i_0a, simp11_0[0:0], simp11_0[1:1]);
endmodule

// tkj32m32_0 TeakJ [Many [32,0],One 32]
module tkj32m32_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_0r1[24:24]);
  BUFF I57 (joint_0[25:25], i_0r1[25:25]);
  BUFF I58 (joint_0[26:26], i_0r1[26:26]);
  BUFF I59 (joint_0[27:27], i_0r1[27:27]);
  BUFF I60 (joint_0[28:28], i_0r1[28:28]);
  BUFF I61 (joint_0[29:29], i_0r1[29:29]);
  BUFF I62 (joint_0[30:30], i_0r1[30:30]);
  BUFF I63 (joint_0[31:31], i_0r1[31:31]);
  BUFF I64 (icomplete_0, i_1r);
  C2 I65 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I66 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I67 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I68 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I69 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I70 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I71 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I72 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I73 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I74 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I75 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I76 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I77 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I78 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I79 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I80 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I81 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I82 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I83 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I84 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I85 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I86 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I87 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I88 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I89 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I90 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I91 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I92 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I93 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I94 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I95 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I96 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I97 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I98 (o_0r1[1:1], joint_0[1:1]);
  BUFF I99 (o_0r1[2:2], joint_0[2:2]);
  BUFF I100 (o_0r1[3:3], joint_0[3:3]);
  BUFF I101 (o_0r1[4:4], joint_0[4:4]);
  BUFF I102 (o_0r1[5:5], joint_0[5:5]);
  BUFF I103 (o_0r1[6:6], joint_0[6:6]);
  BUFF I104 (o_0r1[7:7], joint_0[7:7]);
  BUFF I105 (o_0r1[8:8], joint_0[8:8]);
  BUFF I106 (o_0r1[9:9], joint_0[9:9]);
  BUFF I107 (o_0r1[10:10], joint_0[10:10]);
  BUFF I108 (o_0r1[11:11], joint_0[11:11]);
  BUFF I109 (o_0r1[12:12], joint_0[12:12]);
  BUFF I110 (o_0r1[13:13], joint_0[13:13]);
  BUFF I111 (o_0r1[14:14], joint_0[14:14]);
  BUFF I112 (o_0r1[15:15], joint_0[15:15]);
  BUFF I113 (o_0r1[16:16], joint_0[16:16]);
  BUFF I114 (o_0r1[17:17], joint_0[17:17]);
  BUFF I115 (o_0r1[18:18], joint_0[18:18]);
  BUFF I116 (o_0r1[19:19], joint_0[19:19]);
  BUFF I117 (o_0r1[20:20], joint_0[20:20]);
  BUFF I118 (o_0r1[21:21], joint_0[21:21]);
  BUFF I119 (o_0r1[22:22], joint_0[22:22]);
  BUFF I120 (o_0r1[23:23], joint_0[23:23]);
  BUFF I121 (o_0r1[24:24], joint_0[24:24]);
  BUFF I122 (o_0r1[25:25], joint_0[25:25]);
  BUFF I123 (o_0r1[26:26], joint_0[26:26]);
  BUFF I124 (o_0r1[27:27], joint_0[27:27]);
  BUFF I125 (o_0r1[28:28], joint_0[28:28]);
  BUFF I126 (o_0r1[29:29], joint_0[29:29]);
  BUFF I127 (o_0r1[30:30], joint_0[30:30]);
  BUFF I128 (o_0r1[31:31], joint_0[31:31]);
  BUFF I129 (i_0a, o_0a);
  BUFF I130 (i_1a, o_0a);
endmodule

// tkj35m32_3 TeakJ [Many [32,3],One 35]
module tkj35m32_3 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [34:0] o_0r0;
  output [34:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [34:0] joinf_0;
  wire [34:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joinf_0[34:34], i_1r0[2:2]);
  BUFF I35 (joint_0[0:0], i_0r1[0:0]);
  BUFF I36 (joint_0[1:1], i_0r1[1:1]);
  BUFF I37 (joint_0[2:2], i_0r1[2:2]);
  BUFF I38 (joint_0[3:3], i_0r1[3:3]);
  BUFF I39 (joint_0[4:4], i_0r1[4:4]);
  BUFF I40 (joint_0[5:5], i_0r1[5:5]);
  BUFF I41 (joint_0[6:6], i_0r1[6:6]);
  BUFF I42 (joint_0[7:7], i_0r1[7:7]);
  BUFF I43 (joint_0[8:8], i_0r1[8:8]);
  BUFF I44 (joint_0[9:9], i_0r1[9:9]);
  BUFF I45 (joint_0[10:10], i_0r1[10:10]);
  BUFF I46 (joint_0[11:11], i_0r1[11:11]);
  BUFF I47 (joint_0[12:12], i_0r1[12:12]);
  BUFF I48 (joint_0[13:13], i_0r1[13:13]);
  BUFF I49 (joint_0[14:14], i_0r1[14:14]);
  BUFF I50 (joint_0[15:15], i_0r1[15:15]);
  BUFF I51 (joint_0[16:16], i_0r1[16:16]);
  BUFF I52 (joint_0[17:17], i_0r1[17:17]);
  BUFF I53 (joint_0[18:18], i_0r1[18:18]);
  BUFF I54 (joint_0[19:19], i_0r1[19:19]);
  BUFF I55 (joint_0[20:20], i_0r1[20:20]);
  BUFF I56 (joint_0[21:21], i_0r1[21:21]);
  BUFF I57 (joint_0[22:22], i_0r1[22:22]);
  BUFF I58 (joint_0[23:23], i_0r1[23:23]);
  BUFF I59 (joint_0[24:24], i_0r1[24:24]);
  BUFF I60 (joint_0[25:25], i_0r1[25:25]);
  BUFF I61 (joint_0[26:26], i_0r1[26:26]);
  BUFF I62 (joint_0[27:27], i_0r1[27:27]);
  BUFF I63 (joint_0[28:28], i_0r1[28:28]);
  BUFF I64 (joint_0[29:29], i_0r1[29:29]);
  BUFF I65 (joint_0[30:30], i_0r1[30:30]);
  BUFF I66 (joint_0[31:31], i_0r1[31:31]);
  BUFF I67 (joint_0[32:32], i_1r1[0:0]);
  BUFF I68 (joint_0[33:33], i_1r1[1:1]);
  BUFF I69 (joint_0[34:34], i_1r1[2:2]);
  OR2 I70 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I71 (icomplete_0, dcomplete_0);
  C2 I72 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I73 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I74 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I75 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I76 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I77 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I78 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I79 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I80 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I81 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I82 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I83 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I84 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I85 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I86 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I87 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I88 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I89 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I90 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I91 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I92 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I93 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I94 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I95 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I96 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I97 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I98 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I99 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I100 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I101 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I102 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I103 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I104 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I105 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I106 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I107 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I108 (o_0r1[1:1], joint_0[1:1]);
  BUFF I109 (o_0r1[2:2], joint_0[2:2]);
  BUFF I110 (o_0r1[3:3], joint_0[3:3]);
  BUFF I111 (o_0r1[4:4], joint_0[4:4]);
  BUFF I112 (o_0r1[5:5], joint_0[5:5]);
  BUFF I113 (o_0r1[6:6], joint_0[6:6]);
  BUFF I114 (o_0r1[7:7], joint_0[7:7]);
  BUFF I115 (o_0r1[8:8], joint_0[8:8]);
  BUFF I116 (o_0r1[9:9], joint_0[9:9]);
  BUFF I117 (o_0r1[10:10], joint_0[10:10]);
  BUFF I118 (o_0r1[11:11], joint_0[11:11]);
  BUFF I119 (o_0r1[12:12], joint_0[12:12]);
  BUFF I120 (o_0r1[13:13], joint_0[13:13]);
  BUFF I121 (o_0r1[14:14], joint_0[14:14]);
  BUFF I122 (o_0r1[15:15], joint_0[15:15]);
  BUFF I123 (o_0r1[16:16], joint_0[16:16]);
  BUFF I124 (o_0r1[17:17], joint_0[17:17]);
  BUFF I125 (o_0r1[18:18], joint_0[18:18]);
  BUFF I126 (o_0r1[19:19], joint_0[19:19]);
  BUFF I127 (o_0r1[20:20], joint_0[20:20]);
  BUFF I128 (o_0r1[21:21], joint_0[21:21]);
  BUFF I129 (o_0r1[22:22], joint_0[22:22]);
  BUFF I130 (o_0r1[23:23], joint_0[23:23]);
  BUFF I131 (o_0r1[24:24], joint_0[24:24]);
  BUFF I132 (o_0r1[25:25], joint_0[25:25]);
  BUFF I133 (o_0r1[26:26], joint_0[26:26]);
  BUFF I134 (o_0r1[27:27], joint_0[27:27]);
  BUFF I135 (o_0r1[28:28], joint_0[28:28]);
  BUFF I136 (o_0r1[29:29], joint_0[29:29]);
  BUFF I137 (o_0r1[30:30], joint_0[30:30]);
  BUFF I138 (o_0r1[31:31], joint_0[31:31]);
  BUFF I139 (o_0r1[32:32], joint_0[32:32]);
  BUFF I140 (o_0r1[33:33], joint_0[33:33]);
  BUFF I141 (o_0r1[34:34], joint_0[34:34]);
  BUFF I142 (i_0a, o_0a);
  BUFF I143 (i_1a, o_0a);
endmodule

// tks35_o32w3_1o0w32_2o0w32_4o0w32 TeakS (32+:3) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0)] [One 35,M
//   any [32,32,32]]
module tks35_o32w3_1o0w32_2o0w32_4o0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, reset);
  input [34:0] i_0r0;
  input [34:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  output [31:0] o_2r0;
  output [31:0] o_2r1;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [34:0] comp_0;
  wire [11:0] simp561_0;
  wire [3:0] simp562_0;
  wire [1:0] simp563_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[32:32], i_0r0[33:33], i_0r0[34:34]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[32:32], i_0r0[33:33], i_0r1[34:34]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I11 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I12 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I13 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I14 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I15 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I16 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I17 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I18 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I19 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I20 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I21 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I22 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I23 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I24 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I25 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I26 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I27 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I28 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I29 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I30 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I31 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I32 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I33 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I34 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I35 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I36 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I37 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I38 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I39 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I40 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I41 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I42 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I43 (comp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  C3 I44 (simp561_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I45 (simp561_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I46 (simp561_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I47 (simp561_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I48 (simp561_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I49 (simp561_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I50 (simp561_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I51 (simp561_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I52 (simp561_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I53 (simp561_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I54 (simp561_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  C2 I55 (simp561_0[11:11], comp_0[33:33], comp_0[34:34]);
  C3 I56 (simp562_0[0:0], simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  C3 I57 (simp562_0[1:1], simp561_0[3:3], simp561_0[4:4], simp561_0[5:5]);
  C3 I58 (simp562_0[2:2], simp561_0[6:6], simp561_0[7:7], simp561_0[8:8]);
  C3 I59 (simp562_0[3:3], simp561_0[9:9], simp561_0[10:10], simp561_0[11:11]);
  C3 I60 (simp563_0[0:0], simp562_0[0:0], simp562_0[1:1], simp562_0[2:2]);
  BUFF I61 (simp563_0[1:1], simp562_0[3:3]);
  C2 I62 (icomplete_0, simp563_0[0:0], simp563_0[1:1]);
  C2 I63 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I64 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I65 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I66 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I67 (o_0r0[4:4], i_0r0[4:4], gsel_0);
  C2 I68 (o_0r0[5:5], i_0r0[5:5], gsel_0);
  C2 I69 (o_0r0[6:6], i_0r0[6:6], gsel_0);
  C2 I70 (o_0r0[7:7], i_0r0[7:7], gsel_0);
  C2 I71 (o_0r0[8:8], i_0r0[8:8], gsel_0);
  C2 I72 (o_0r0[9:9], i_0r0[9:9], gsel_0);
  C2 I73 (o_0r0[10:10], i_0r0[10:10], gsel_0);
  C2 I74 (o_0r0[11:11], i_0r0[11:11], gsel_0);
  C2 I75 (o_0r0[12:12], i_0r0[12:12], gsel_0);
  C2 I76 (o_0r0[13:13], i_0r0[13:13], gsel_0);
  C2 I77 (o_0r0[14:14], i_0r0[14:14], gsel_0);
  C2 I78 (o_0r0[15:15], i_0r0[15:15], gsel_0);
  C2 I79 (o_0r0[16:16], i_0r0[16:16], gsel_0);
  C2 I80 (o_0r0[17:17], i_0r0[17:17], gsel_0);
  C2 I81 (o_0r0[18:18], i_0r0[18:18], gsel_0);
  C2 I82 (o_0r0[19:19], i_0r0[19:19], gsel_0);
  C2 I83 (o_0r0[20:20], i_0r0[20:20], gsel_0);
  C2 I84 (o_0r0[21:21], i_0r0[21:21], gsel_0);
  C2 I85 (o_0r0[22:22], i_0r0[22:22], gsel_0);
  C2 I86 (o_0r0[23:23], i_0r0[23:23], gsel_0);
  C2 I87 (o_0r0[24:24], i_0r0[24:24], gsel_0);
  C2 I88 (o_0r0[25:25], i_0r0[25:25], gsel_0);
  C2 I89 (o_0r0[26:26], i_0r0[26:26], gsel_0);
  C2 I90 (o_0r0[27:27], i_0r0[27:27], gsel_0);
  C2 I91 (o_0r0[28:28], i_0r0[28:28], gsel_0);
  C2 I92 (o_0r0[29:29], i_0r0[29:29], gsel_0);
  C2 I93 (o_0r0[30:30], i_0r0[30:30], gsel_0);
  C2 I94 (o_0r0[31:31], i_0r0[31:31], gsel_0);
  C2 I95 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I96 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I97 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I98 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I99 (o_1r0[4:4], i_0r0[4:4], gsel_1);
  C2 I100 (o_1r0[5:5], i_0r0[5:5], gsel_1);
  C2 I101 (o_1r0[6:6], i_0r0[6:6], gsel_1);
  C2 I102 (o_1r0[7:7], i_0r0[7:7], gsel_1);
  C2 I103 (o_1r0[8:8], i_0r0[8:8], gsel_1);
  C2 I104 (o_1r0[9:9], i_0r0[9:9], gsel_1);
  C2 I105 (o_1r0[10:10], i_0r0[10:10], gsel_1);
  C2 I106 (o_1r0[11:11], i_0r0[11:11], gsel_1);
  C2 I107 (o_1r0[12:12], i_0r0[12:12], gsel_1);
  C2 I108 (o_1r0[13:13], i_0r0[13:13], gsel_1);
  C2 I109 (o_1r0[14:14], i_0r0[14:14], gsel_1);
  C2 I110 (o_1r0[15:15], i_0r0[15:15], gsel_1);
  C2 I111 (o_1r0[16:16], i_0r0[16:16], gsel_1);
  C2 I112 (o_1r0[17:17], i_0r0[17:17], gsel_1);
  C2 I113 (o_1r0[18:18], i_0r0[18:18], gsel_1);
  C2 I114 (o_1r0[19:19], i_0r0[19:19], gsel_1);
  C2 I115 (o_1r0[20:20], i_0r0[20:20], gsel_1);
  C2 I116 (o_1r0[21:21], i_0r0[21:21], gsel_1);
  C2 I117 (o_1r0[22:22], i_0r0[22:22], gsel_1);
  C2 I118 (o_1r0[23:23], i_0r0[23:23], gsel_1);
  C2 I119 (o_1r0[24:24], i_0r0[24:24], gsel_1);
  C2 I120 (o_1r0[25:25], i_0r0[25:25], gsel_1);
  C2 I121 (o_1r0[26:26], i_0r0[26:26], gsel_1);
  C2 I122 (o_1r0[27:27], i_0r0[27:27], gsel_1);
  C2 I123 (o_1r0[28:28], i_0r0[28:28], gsel_1);
  C2 I124 (o_1r0[29:29], i_0r0[29:29], gsel_1);
  C2 I125 (o_1r0[30:30], i_0r0[30:30], gsel_1);
  C2 I126 (o_1r0[31:31], i_0r0[31:31], gsel_1);
  C2 I127 (o_2r0[0:0], i_0r0[0:0], gsel_2);
  C2 I128 (o_2r0[1:1], i_0r0[1:1], gsel_2);
  C2 I129 (o_2r0[2:2], i_0r0[2:2], gsel_2);
  C2 I130 (o_2r0[3:3], i_0r0[3:3], gsel_2);
  C2 I131 (o_2r0[4:4], i_0r0[4:4], gsel_2);
  C2 I132 (o_2r0[5:5], i_0r0[5:5], gsel_2);
  C2 I133 (o_2r0[6:6], i_0r0[6:6], gsel_2);
  C2 I134 (o_2r0[7:7], i_0r0[7:7], gsel_2);
  C2 I135 (o_2r0[8:8], i_0r0[8:8], gsel_2);
  C2 I136 (o_2r0[9:9], i_0r0[9:9], gsel_2);
  C2 I137 (o_2r0[10:10], i_0r0[10:10], gsel_2);
  C2 I138 (o_2r0[11:11], i_0r0[11:11], gsel_2);
  C2 I139 (o_2r0[12:12], i_0r0[12:12], gsel_2);
  C2 I140 (o_2r0[13:13], i_0r0[13:13], gsel_2);
  C2 I141 (o_2r0[14:14], i_0r0[14:14], gsel_2);
  C2 I142 (o_2r0[15:15], i_0r0[15:15], gsel_2);
  C2 I143 (o_2r0[16:16], i_0r0[16:16], gsel_2);
  C2 I144 (o_2r0[17:17], i_0r0[17:17], gsel_2);
  C2 I145 (o_2r0[18:18], i_0r0[18:18], gsel_2);
  C2 I146 (o_2r0[19:19], i_0r0[19:19], gsel_2);
  C2 I147 (o_2r0[20:20], i_0r0[20:20], gsel_2);
  C2 I148 (o_2r0[21:21], i_0r0[21:21], gsel_2);
  C2 I149 (o_2r0[22:22], i_0r0[22:22], gsel_2);
  C2 I150 (o_2r0[23:23], i_0r0[23:23], gsel_2);
  C2 I151 (o_2r0[24:24], i_0r0[24:24], gsel_2);
  C2 I152 (o_2r0[25:25], i_0r0[25:25], gsel_2);
  C2 I153 (o_2r0[26:26], i_0r0[26:26], gsel_2);
  C2 I154 (o_2r0[27:27], i_0r0[27:27], gsel_2);
  C2 I155 (o_2r0[28:28], i_0r0[28:28], gsel_2);
  C2 I156 (o_2r0[29:29], i_0r0[29:29], gsel_2);
  C2 I157 (o_2r0[30:30], i_0r0[30:30], gsel_2);
  C2 I158 (o_2r0[31:31], i_0r0[31:31], gsel_2);
  C2 I159 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I160 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I161 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I162 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I163 (o_0r1[4:4], i_0r1[4:4], gsel_0);
  C2 I164 (o_0r1[5:5], i_0r1[5:5], gsel_0);
  C2 I165 (o_0r1[6:6], i_0r1[6:6], gsel_0);
  C2 I166 (o_0r1[7:7], i_0r1[7:7], gsel_0);
  C2 I167 (o_0r1[8:8], i_0r1[8:8], gsel_0);
  C2 I168 (o_0r1[9:9], i_0r1[9:9], gsel_0);
  C2 I169 (o_0r1[10:10], i_0r1[10:10], gsel_0);
  C2 I170 (o_0r1[11:11], i_0r1[11:11], gsel_0);
  C2 I171 (o_0r1[12:12], i_0r1[12:12], gsel_0);
  C2 I172 (o_0r1[13:13], i_0r1[13:13], gsel_0);
  C2 I173 (o_0r1[14:14], i_0r1[14:14], gsel_0);
  C2 I174 (o_0r1[15:15], i_0r1[15:15], gsel_0);
  C2 I175 (o_0r1[16:16], i_0r1[16:16], gsel_0);
  C2 I176 (o_0r1[17:17], i_0r1[17:17], gsel_0);
  C2 I177 (o_0r1[18:18], i_0r1[18:18], gsel_0);
  C2 I178 (o_0r1[19:19], i_0r1[19:19], gsel_0);
  C2 I179 (o_0r1[20:20], i_0r1[20:20], gsel_0);
  C2 I180 (o_0r1[21:21], i_0r1[21:21], gsel_0);
  C2 I181 (o_0r1[22:22], i_0r1[22:22], gsel_0);
  C2 I182 (o_0r1[23:23], i_0r1[23:23], gsel_0);
  C2 I183 (o_0r1[24:24], i_0r1[24:24], gsel_0);
  C2 I184 (o_0r1[25:25], i_0r1[25:25], gsel_0);
  C2 I185 (o_0r1[26:26], i_0r1[26:26], gsel_0);
  C2 I186 (o_0r1[27:27], i_0r1[27:27], gsel_0);
  C2 I187 (o_0r1[28:28], i_0r1[28:28], gsel_0);
  C2 I188 (o_0r1[29:29], i_0r1[29:29], gsel_0);
  C2 I189 (o_0r1[30:30], i_0r1[30:30], gsel_0);
  C2 I190 (o_0r1[31:31], i_0r1[31:31], gsel_0);
  C2 I191 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I192 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I193 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I194 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I195 (o_1r1[4:4], i_0r1[4:4], gsel_1);
  C2 I196 (o_1r1[5:5], i_0r1[5:5], gsel_1);
  C2 I197 (o_1r1[6:6], i_0r1[6:6], gsel_1);
  C2 I198 (o_1r1[7:7], i_0r1[7:7], gsel_1);
  C2 I199 (o_1r1[8:8], i_0r1[8:8], gsel_1);
  C2 I200 (o_1r1[9:9], i_0r1[9:9], gsel_1);
  C2 I201 (o_1r1[10:10], i_0r1[10:10], gsel_1);
  C2 I202 (o_1r1[11:11], i_0r1[11:11], gsel_1);
  C2 I203 (o_1r1[12:12], i_0r1[12:12], gsel_1);
  C2 I204 (o_1r1[13:13], i_0r1[13:13], gsel_1);
  C2 I205 (o_1r1[14:14], i_0r1[14:14], gsel_1);
  C2 I206 (o_1r1[15:15], i_0r1[15:15], gsel_1);
  C2 I207 (o_1r1[16:16], i_0r1[16:16], gsel_1);
  C2 I208 (o_1r1[17:17], i_0r1[17:17], gsel_1);
  C2 I209 (o_1r1[18:18], i_0r1[18:18], gsel_1);
  C2 I210 (o_1r1[19:19], i_0r1[19:19], gsel_1);
  C2 I211 (o_1r1[20:20], i_0r1[20:20], gsel_1);
  C2 I212 (o_1r1[21:21], i_0r1[21:21], gsel_1);
  C2 I213 (o_1r1[22:22], i_0r1[22:22], gsel_1);
  C2 I214 (o_1r1[23:23], i_0r1[23:23], gsel_1);
  C2 I215 (o_1r1[24:24], i_0r1[24:24], gsel_1);
  C2 I216 (o_1r1[25:25], i_0r1[25:25], gsel_1);
  C2 I217 (o_1r1[26:26], i_0r1[26:26], gsel_1);
  C2 I218 (o_1r1[27:27], i_0r1[27:27], gsel_1);
  C2 I219 (o_1r1[28:28], i_0r1[28:28], gsel_1);
  C2 I220 (o_1r1[29:29], i_0r1[29:29], gsel_1);
  C2 I221 (o_1r1[30:30], i_0r1[30:30], gsel_1);
  C2 I222 (o_1r1[31:31], i_0r1[31:31], gsel_1);
  C2 I223 (o_2r1[0:0], i_0r1[0:0], gsel_2);
  C2 I224 (o_2r1[1:1], i_0r1[1:1], gsel_2);
  C2 I225 (o_2r1[2:2], i_0r1[2:2], gsel_2);
  C2 I226 (o_2r1[3:3], i_0r1[3:3], gsel_2);
  C2 I227 (o_2r1[4:4], i_0r1[4:4], gsel_2);
  C2 I228 (o_2r1[5:5], i_0r1[5:5], gsel_2);
  C2 I229 (o_2r1[6:6], i_0r1[6:6], gsel_2);
  C2 I230 (o_2r1[7:7], i_0r1[7:7], gsel_2);
  C2 I231 (o_2r1[8:8], i_0r1[8:8], gsel_2);
  C2 I232 (o_2r1[9:9], i_0r1[9:9], gsel_2);
  C2 I233 (o_2r1[10:10], i_0r1[10:10], gsel_2);
  C2 I234 (o_2r1[11:11], i_0r1[11:11], gsel_2);
  C2 I235 (o_2r1[12:12], i_0r1[12:12], gsel_2);
  C2 I236 (o_2r1[13:13], i_0r1[13:13], gsel_2);
  C2 I237 (o_2r1[14:14], i_0r1[14:14], gsel_2);
  C2 I238 (o_2r1[15:15], i_0r1[15:15], gsel_2);
  C2 I239 (o_2r1[16:16], i_0r1[16:16], gsel_2);
  C2 I240 (o_2r1[17:17], i_0r1[17:17], gsel_2);
  C2 I241 (o_2r1[18:18], i_0r1[18:18], gsel_2);
  C2 I242 (o_2r1[19:19], i_0r1[19:19], gsel_2);
  C2 I243 (o_2r1[20:20], i_0r1[20:20], gsel_2);
  C2 I244 (o_2r1[21:21], i_0r1[21:21], gsel_2);
  C2 I245 (o_2r1[22:22], i_0r1[22:22], gsel_2);
  C2 I246 (o_2r1[23:23], i_0r1[23:23], gsel_2);
  C2 I247 (o_2r1[24:24], i_0r1[24:24], gsel_2);
  C2 I248 (o_2r1[25:25], i_0r1[25:25], gsel_2);
  C2 I249 (o_2r1[26:26], i_0r1[26:26], gsel_2);
  C2 I250 (o_2r1[27:27], i_0r1[27:27], gsel_2);
  C2 I251 (o_2r1[28:28], i_0r1[28:28], gsel_2);
  C2 I252 (o_2r1[29:29], i_0r1[29:29], gsel_2);
  C2 I253 (o_2r1[30:30], i_0r1[30:30], gsel_2);
  C2 I254 (o_2r1[31:31], i_0r1[31:31], gsel_2);
  OR3 I255 (oack_0, o_0a, o_1a, o_2a);
  C2 I256 (i_0a, oack_0, icomplete_0);
endmodule

// tkvxV32_wo0w32_ro0w32 TeakV "xV" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvxV32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w32o31w1 TeakV "i" 32 [] [0] [0,0,31] [Many [32],Many [0],Many [0,0,0],Many [3
//   2,32,1]]
module tkvi32_wo0w32_ro0w32o0w32o31w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp5381_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0, df_0[31:31], rg_2r);
  AND2 I489 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I490 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I491 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I492 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I493 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I494 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I495 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I496 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I497 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I498 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I499 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I500 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I501 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I502 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I503 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I504 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I505 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I506 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I507 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I508 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I509 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I510 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I511 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I512 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I513 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I514 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I515 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I516 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I517 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I518 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I519 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I520 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I521 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I522 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I523 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I524 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I525 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I526 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I527 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I528 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I529 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I530 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I531 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I532 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I533 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I534 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I535 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I536 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I537 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I538 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I539 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I540 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I541 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I542 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I543 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I544 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I545 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I546 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I547 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I548 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I549 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I550 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I551 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I552 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I553 (rd_2r1, dt_0[31:31], rg_2r);
  NOR3 I554 (simp5381_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I555 (simp5381_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I556 (anyread_0, simp5381_0[0:0], simp5381_0[1:1]);
  BUFF I557 (wg_0a, wd_0a);
  BUFF I558 (rg_0a, rd_0a);
  BUFF I559 (rg_1a, rd_1a);
  BUFF I560 (rg_2a, rd_2a);
endmodule

// tkvaV32_wo0w32_ro0w32o0w32 TeakV "aV" 32 [] [0] [0,0] [Many [32],Many [0],Many [0,0],Many [32,32]]
module tkvaV32_wo0w32_ro0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp5361_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I489 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I490 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I491 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I492 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I493 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I494 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I495 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I496 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I497 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I498 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I499 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I500 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I501 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I502 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I503 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I504 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I505 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I506 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I507 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I508 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I509 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I510 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I511 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I512 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I513 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I514 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I515 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I516 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I517 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I518 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I519 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I520 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I521 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I522 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I523 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I524 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I525 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I526 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I527 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I528 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I529 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I530 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I531 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I532 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I533 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I534 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I535 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I536 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I537 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I538 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I539 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I540 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I541 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I542 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I543 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I544 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I545 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I546 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I547 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I548 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I549 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I550 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I551 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  NOR3 I552 (simp5361_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I553 (simp5361_0[1:1], rg_1a);
  NAND2 I554 (anyread_0, simp5361_0[0:0], simp5361_0[1:1]);
  BUFF I555 (wg_0a, wd_0a);
  BUFF I556 (rg_0a, rd_0a);
  BUFF I557 (rg_1a, rd_1a);
endmodule

// tkj34m32_2 TeakJ [Many [32,2],One 34]
module tkj34m32_2 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [33:0] o_0r0;
  output [33:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [33:0] joinf_0;
  wire [33:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joint_0[0:0], i_0r1[0:0]);
  BUFF I35 (joint_0[1:1], i_0r1[1:1]);
  BUFF I36 (joint_0[2:2], i_0r1[2:2]);
  BUFF I37 (joint_0[3:3], i_0r1[3:3]);
  BUFF I38 (joint_0[4:4], i_0r1[4:4]);
  BUFF I39 (joint_0[5:5], i_0r1[5:5]);
  BUFF I40 (joint_0[6:6], i_0r1[6:6]);
  BUFF I41 (joint_0[7:7], i_0r1[7:7]);
  BUFF I42 (joint_0[8:8], i_0r1[8:8]);
  BUFF I43 (joint_0[9:9], i_0r1[9:9]);
  BUFF I44 (joint_0[10:10], i_0r1[10:10]);
  BUFF I45 (joint_0[11:11], i_0r1[11:11]);
  BUFF I46 (joint_0[12:12], i_0r1[12:12]);
  BUFF I47 (joint_0[13:13], i_0r1[13:13]);
  BUFF I48 (joint_0[14:14], i_0r1[14:14]);
  BUFF I49 (joint_0[15:15], i_0r1[15:15]);
  BUFF I50 (joint_0[16:16], i_0r1[16:16]);
  BUFF I51 (joint_0[17:17], i_0r1[17:17]);
  BUFF I52 (joint_0[18:18], i_0r1[18:18]);
  BUFF I53 (joint_0[19:19], i_0r1[19:19]);
  BUFF I54 (joint_0[20:20], i_0r1[20:20]);
  BUFF I55 (joint_0[21:21], i_0r1[21:21]);
  BUFF I56 (joint_0[22:22], i_0r1[22:22]);
  BUFF I57 (joint_0[23:23], i_0r1[23:23]);
  BUFF I58 (joint_0[24:24], i_0r1[24:24]);
  BUFF I59 (joint_0[25:25], i_0r1[25:25]);
  BUFF I60 (joint_0[26:26], i_0r1[26:26]);
  BUFF I61 (joint_0[27:27], i_0r1[27:27]);
  BUFF I62 (joint_0[28:28], i_0r1[28:28]);
  BUFF I63 (joint_0[29:29], i_0r1[29:29]);
  BUFF I64 (joint_0[30:30], i_0r1[30:30]);
  BUFF I65 (joint_0[31:31], i_0r1[31:31]);
  BUFF I66 (joint_0[32:32], i_1r1[0:0]);
  BUFF I67 (joint_0[33:33], i_1r1[1:1]);
  OR2 I68 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I69 (icomplete_0, dcomplete_0);
  C2 I70 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I71 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I72 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I73 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I74 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I75 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I76 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I77 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I78 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I79 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I80 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I81 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I82 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I83 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I84 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I85 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I86 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I87 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I88 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I89 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I90 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I91 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I92 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I93 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I94 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I95 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I96 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I97 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I98 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I99 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I100 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I101 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I102 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I103 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I104 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I105 (o_0r1[1:1], joint_0[1:1]);
  BUFF I106 (o_0r1[2:2], joint_0[2:2]);
  BUFF I107 (o_0r1[3:3], joint_0[3:3]);
  BUFF I108 (o_0r1[4:4], joint_0[4:4]);
  BUFF I109 (o_0r1[5:5], joint_0[5:5]);
  BUFF I110 (o_0r1[6:6], joint_0[6:6]);
  BUFF I111 (o_0r1[7:7], joint_0[7:7]);
  BUFF I112 (o_0r1[8:8], joint_0[8:8]);
  BUFF I113 (o_0r1[9:9], joint_0[9:9]);
  BUFF I114 (o_0r1[10:10], joint_0[10:10]);
  BUFF I115 (o_0r1[11:11], joint_0[11:11]);
  BUFF I116 (o_0r1[12:12], joint_0[12:12]);
  BUFF I117 (o_0r1[13:13], joint_0[13:13]);
  BUFF I118 (o_0r1[14:14], joint_0[14:14]);
  BUFF I119 (o_0r1[15:15], joint_0[15:15]);
  BUFF I120 (o_0r1[16:16], joint_0[16:16]);
  BUFF I121 (o_0r1[17:17], joint_0[17:17]);
  BUFF I122 (o_0r1[18:18], joint_0[18:18]);
  BUFF I123 (o_0r1[19:19], joint_0[19:19]);
  BUFF I124 (o_0r1[20:20], joint_0[20:20]);
  BUFF I125 (o_0r1[21:21], joint_0[21:21]);
  BUFF I126 (o_0r1[22:22], joint_0[22:22]);
  BUFF I127 (o_0r1[23:23], joint_0[23:23]);
  BUFF I128 (o_0r1[24:24], joint_0[24:24]);
  BUFF I129 (o_0r1[25:25], joint_0[25:25]);
  BUFF I130 (o_0r1[26:26], joint_0[26:26]);
  BUFF I131 (o_0r1[27:27], joint_0[27:27]);
  BUFF I132 (o_0r1[28:28], joint_0[28:28]);
  BUFF I133 (o_0r1[29:29], joint_0[29:29]);
  BUFF I134 (o_0r1[30:30], joint_0[30:30]);
  BUFF I135 (o_0r1[31:31], joint_0[31:31]);
  BUFF I136 (o_0r1[32:32], joint_0[32:32]);
  BUFF I137 (o_0r1[33:33], joint_0[33:33]);
  BUFF I138 (i_0a, o_0a);
  BUFF I139 (i_1a, o_0a);
endmodule

// tks34_o32w2_1o0w32_2o0w32 TeakS (32+:2) [([Imp 1 0],0),([Imp 2 0],0)] [One 34,Many [32,32]]
module tks34_o32w2_1o0w32_2o0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [33:0] i_0r0;
  input [33:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire [33:0] comp_0;
  wire [11:0] simp491_0;
  wire [3:0] simp492_0;
  wire [1:0] simp493_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[32:32], i_0r0[33:33]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r0[32:32], i_0r1[33:33]);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I7 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I8 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I9 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I10 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I11 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I12 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I13 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I14 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I15 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I16 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I17 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I18 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I19 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I20 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I21 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I22 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I23 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I24 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I25 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I26 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I27 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I28 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I29 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I30 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I31 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I32 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I33 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I34 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I35 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I36 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I37 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I38 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I39 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  C3 I40 (simp491_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I41 (simp491_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I42 (simp491_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I43 (simp491_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I44 (simp491_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I45 (simp491_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I46 (simp491_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I47 (simp491_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I48 (simp491_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I49 (simp491_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I50 (simp491_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  BUFF I51 (simp491_0[11:11], comp_0[33:33]);
  C3 I52 (simp492_0[0:0], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  C3 I53 (simp492_0[1:1], simp491_0[3:3], simp491_0[4:4], simp491_0[5:5]);
  C3 I54 (simp492_0[2:2], simp491_0[6:6], simp491_0[7:7], simp491_0[8:8]);
  C3 I55 (simp492_0[3:3], simp491_0[9:9], simp491_0[10:10], simp491_0[11:11]);
  C3 I56 (simp493_0[0:0], simp492_0[0:0], simp492_0[1:1], simp492_0[2:2]);
  BUFF I57 (simp493_0[1:1], simp492_0[3:3]);
  C2 I58 (icomplete_0, simp493_0[0:0], simp493_0[1:1]);
  C2 I59 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I60 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I61 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I62 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I63 (o_0r0[4:4], i_0r0[4:4], gsel_0);
  C2 I64 (o_0r0[5:5], i_0r0[5:5], gsel_0);
  C2 I65 (o_0r0[6:6], i_0r0[6:6], gsel_0);
  C2 I66 (o_0r0[7:7], i_0r0[7:7], gsel_0);
  C2 I67 (o_0r0[8:8], i_0r0[8:8], gsel_0);
  C2 I68 (o_0r0[9:9], i_0r0[9:9], gsel_0);
  C2 I69 (o_0r0[10:10], i_0r0[10:10], gsel_0);
  C2 I70 (o_0r0[11:11], i_0r0[11:11], gsel_0);
  C2 I71 (o_0r0[12:12], i_0r0[12:12], gsel_0);
  C2 I72 (o_0r0[13:13], i_0r0[13:13], gsel_0);
  C2 I73 (o_0r0[14:14], i_0r0[14:14], gsel_0);
  C2 I74 (o_0r0[15:15], i_0r0[15:15], gsel_0);
  C2 I75 (o_0r0[16:16], i_0r0[16:16], gsel_0);
  C2 I76 (o_0r0[17:17], i_0r0[17:17], gsel_0);
  C2 I77 (o_0r0[18:18], i_0r0[18:18], gsel_0);
  C2 I78 (o_0r0[19:19], i_0r0[19:19], gsel_0);
  C2 I79 (o_0r0[20:20], i_0r0[20:20], gsel_0);
  C2 I80 (o_0r0[21:21], i_0r0[21:21], gsel_0);
  C2 I81 (o_0r0[22:22], i_0r0[22:22], gsel_0);
  C2 I82 (o_0r0[23:23], i_0r0[23:23], gsel_0);
  C2 I83 (o_0r0[24:24], i_0r0[24:24], gsel_0);
  C2 I84 (o_0r0[25:25], i_0r0[25:25], gsel_0);
  C2 I85 (o_0r0[26:26], i_0r0[26:26], gsel_0);
  C2 I86 (o_0r0[27:27], i_0r0[27:27], gsel_0);
  C2 I87 (o_0r0[28:28], i_0r0[28:28], gsel_0);
  C2 I88 (o_0r0[29:29], i_0r0[29:29], gsel_0);
  C2 I89 (o_0r0[30:30], i_0r0[30:30], gsel_0);
  C2 I90 (o_0r0[31:31], i_0r0[31:31], gsel_0);
  C2 I91 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I92 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I93 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I94 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I95 (o_1r0[4:4], i_0r0[4:4], gsel_1);
  C2 I96 (o_1r0[5:5], i_0r0[5:5], gsel_1);
  C2 I97 (o_1r0[6:6], i_0r0[6:6], gsel_1);
  C2 I98 (o_1r0[7:7], i_0r0[7:7], gsel_1);
  C2 I99 (o_1r0[8:8], i_0r0[8:8], gsel_1);
  C2 I100 (o_1r0[9:9], i_0r0[9:9], gsel_1);
  C2 I101 (o_1r0[10:10], i_0r0[10:10], gsel_1);
  C2 I102 (o_1r0[11:11], i_0r0[11:11], gsel_1);
  C2 I103 (o_1r0[12:12], i_0r0[12:12], gsel_1);
  C2 I104 (o_1r0[13:13], i_0r0[13:13], gsel_1);
  C2 I105 (o_1r0[14:14], i_0r0[14:14], gsel_1);
  C2 I106 (o_1r0[15:15], i_0r0[15:15], gsel_1);
  C2 I107 (o_1r0[16:16], i_0r0[16:16], gsel_1);
  C2 I108 (o_1r0[17:17], i_0r0[17:17], gsel_1);
  C2 I109 (o_1r0[18:18], i_0r0[18:18], gsel_1);
  C2 I110 (o_1r0[19:19], i_0r0[19:19], gsel_1);
  C2 I111 (o_1r0[20:20], i_0r0[20:20], gsel_1);
  C2 I112 (o_1r0[21:21], i_0r0[21:21], gsel_1);
  C2 I113 (o_1r0[22:22], i_0r0[22:22], gsel_1);
  C2 I114 (o_1r0[23:23], i_0r0[23:23], gsel_1);
  C2 I115 (o_1r0[24:24], i_0r0[24:24], gsel_1);
  C2 I116 (o_1r0[25:25], i_0r0[25:25], gsel_1);
  C2 I117 (o_1r0[26:26], i_0r0[26:26], gsel_1);
  C2 I118 (o_1r0[27:27], i_0r0[27:27], gsel_1);
  C2 I119 (o_1r0[28:28], i_0r0[28:28], gsel_1);
  C2 I120 (o_1r0[29:29], i_0r0[29:29], gsel_1);
  C2 I121 (o_1r0[30:30], i_0r0[30:30], gsel_1);
  C2 I122 (o_1r0[31:31], i_0r0[31:31], gsel_1);
  C2 I123 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I124 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I125 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I126 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I127 (o_0r1[4:4], i_0r1[4:4], gsel_0);
  C2 I128 (o_0r1[5:5], i_0r1[5:5], gsel_0);
  C2 I129 (o_0r1[6:6], i_0r1[6:6], gsel_0);
  C2 I130 (o_0r1[7:7], i_0r1[7:7], gsel_0);
  C2 I131 (o_0r1[8:8], i_0r1[8:8], gsel_0);
  C2 I132 (o_0r1[9:9], i_0r1[9:9], gsel_0);
  C2 I133 (o_0r1[10:10], i_0r1[10:10], gsel_0);
  C2 I134 (o_0r1[11:11], i_0r1[11:11], gsel_0);
  C2 I135 (o_0r1[12:12], i_0r1[12:12], gsel_0);
  C2 I136 (o_0r1[13:13], i_0r1[13:13], gsel_0);
  C2 I137 (o_0r1[14:14], i_0r1[14:14], gsel_0);
  C2 I138 (o_0r1[15:15], i_0r1[15:15], gsel_0);
  C2 I139 (o_0r1[16:16], i_0r1[16:16], gsel_0);
  C2 I140 (o_0r1[17:17], i_0r1[17:17], gsel_0);
  C2 I141 (o_0r1[18:18], i_0r1[18:18], gsel_0);
  C2 I142 (o_0r1[19:19], i_0r1[19:19], gsel_0);
  C2 I143 (o_0r1[20:20], i_0r1[20:20], gsel_0);
  C2 I144 (o_0r1[21:21], i_0r1[21:21], gsel_0);
  C2 I145 (o_0r1[22:22], i_0r1[22:22], gsel_0);
  C2 I146 (o_0r1[23:23], i_0r1[23:23], gsel_0);
  C2 I147 (o_0r1[24:24], i_0r1[24:24], gsel_0);
  C2 I148 (o_0r1[25:25], i_0r1[25:25], gsel_0);
  C2 I149 (o_0r1[26:26], i_0r1[26:26], gsel_0);
  C2 I150 (o_0r1[27:27], i_0r1[27:27], gsel_0);
  C2 I151 (o_0r1[28:28], i_0r1[28:28], gsel_0);
  C2 I152 (o_0r1[29:29], i_0r1[29:29], gsel_0);
  C2 I153 (o_0r1[30:30], i_0r1[30:30], gsel_0);
  C2 I154 (o_0r1[31:31], i_0r1[31:31], gsel_0);
  C2 I155 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I156 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I157 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I158 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I159 (o_1r1[4:4], i_0r1[4:4], gsel_1);
  C2 I160 (o_1r1[5:5], i_0r1[5:5], gsel_1);
  C2 I161 (o_1r1[6:6], i_0r1[6:6], gsel_1);
  C2 I162 (o_1r1[7:7], i_0r1[7:7], gsel_1);
  C2 I163 (o_1r1[8:8], i_0r1[8:8], gsel_1);
  C2 I164 (o_1r1[9:9], i_0r1[9:9], gsel_1);
  C2 I165 (o_1r1[10:10], i_0r1[10:10], gsel_1);
  C2 I166 (o_1r1[11:11], i_0r1[11:11], gsel_1);
  C2 I167 (o_1r1[12:12], i_0r1[12:12], gsel_1);
  C2 I168 (o_1r1[13:13], i_0r1[13:13], gsel_1);
  C2 I169 (o_1r1[14:14], i_0r1[14:14], gsel_1);
  C2 I170 (o_1r1[15:15], i_0r1[15:15], gsel_1);
  C2 I171 (o_1r1[16:16], i_0r1[16:16], gsel_1);
  C2 I172 (o_1r1[17:17], i_0r1[17:17], gsel_1);
  C2 I173 (o_1r1[18:18], i_0r1[18:18], gsel_1);
  C2 I174 (o_1r1[19:19], i_0r1[19:19], gsel_1);
  C2 I175 (o_1r1[20:20], i_0r1[20:20], gsel_1);
  C2 I176 (o_1r1[21:21], i_0r1[21:21], gsel_1);
  C2 I177 (o_1r1[22:22], i_0r1[22:22], gsel_1);
  C2 I178 (o_1r1[23:23], i_0r1[23:23], gsel_1);
  C2 I179 (o_1r1[24:24], i_0r1[24:24], gsel_1);
  C2 I180 (o_1r1[25:25], i_0r1[25:25], gsel_1);
  C2 I181 (o_1r1[26:26], i_0r1[26:26], gsel_1);
  C2 I182 (o_1r1[27:27], i_0r1[27:27], gsel_1);
  C2 I183 (o_1r1[28:28], i_0r1[28:28], gsel_1);
  C2 I184 (o_1r1[29:29], i_0r1[29:29], gsel_1);
  C2 I185 (o_1r1[30:30], i_0r1[30:30], gsel_1);
  C2 I186 (o_1r1[31:31], i_0r1[31:31], gsel_1);
  OR2 I187 (oack_0, o_0a, o_1a);
  C2 I188 (i_0a, oack_0, icomplete_0);
endmodule

// tki TeakI [One 0,One 0]
module tki (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire nreset_0;
  wire firsthsa_0;
  wire nfirsthsa_0;
  wire firsthsd_0;
  wire noa_0;
  INV I0 (nreset_0, reset);
  INV I1 (nfirsthsa_0, firsthsa_0);
  INV I2 (noa_0, o_0a);
  AO22 I3 (o_0r, nreset_0, nfirsthsa_0, i_0r, firsthsd_0);
  AO22 I4 (firsthsa_0, nreset_0, o_0a, nreset_0, firsthsa_0);
  AO22 I5 (firsthsd_0, firsthsa_0, noa_0, firsthsa_0, firsthsd_0);
  AND2 I6 (i_0a, o_0a, firsthsd_0);
endmodule

// tkj64m32_32_0 TeakJ [Many [32,32,0],One 64]
module tkj64m32_32_0 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input i_2r;
  output i_2a;
  output [63:0] o_0r0;
  output [63:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [63:0] joinf_0;
  wire [63:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joinf_0[34:34], i_1r0[2:2]);
  BUFF I35 (joinf_0[35:35], i_1r0[3:3]);
  BUFF I36 (joinf_0[36:36], i_1r0[4:4]);
  BUFF I37 (joinf_0[37:37], i_1r0[5:5]);
  BUFF I38 (joinf_0[38:38], i_1r0[6:6]);
  BUFF I39 (joinf_0[39:39], i_1r0[7:7]);
  BUFF I40 (joinf_0[40:40], i_1r0[8:8]);
  BUFF I41 (joinf_0[41:41], i_1r0[9:9]);
  BUFF I42 (joinf_0[42:42], i_1r0[10:10]);
  BUFF I43 (joinf_0[43:43], i_1r0[11:11]);
  BUFF I44 (joinf_0[44:44], i_1r0[12:12]);
  BUFF I45 (joinf_0[45:45], i_1r0[13:13]);
  BUFF I46 (joinf_0[46:46], i_1r0[14:14]);
  BUFF I47 (joinf_0[47:47], i_1r0[15:15]);
  BUFF I48 (joinf_0[48:48], i_1r0[16:16]);
  BUFF I49 (joinf_0[49:49], i_1r0[17:17]);
  BUFF I50 (joinf_0[50:50], i_1r0[18:18]);
  BUFF I51 (joinf_0[51:51], i_1r0[19:19]);
  BUFF I52 (joinf_0[52:52], i_1r0[20:20]);
  BUFF I53 (joinf_0[53:53], i_1r0[21:21]);
  BUFF I54 (joinf_0[54:54], i_1r0[22:22]);
  BUFF I55 (joinf_0[55:55], i_1r0[23:23]);
  BUFF I56 (joinf_0[56:56], i_1r0[24:24]);
  BUFF I57 (joinf_0[57:57], i_1r0[25:25]);
  BUFF I58 (joinf_0[58:58], i_1r0[26:26]);
  BUFF I59 (joinf_0[59:59], i_1r0[27:27]);
  BUFF I60 (joinf_0[60:60], i_1r0[28:28]);
  BUFF I61 (joinf_0[61:61], i_1r0[29:29]);
  BUFF I62 (joinf_0[62:62], i_1r0[30:30]);
  BUFF I63 (joinf_0[63:63], i_1r0[31:31]);
  BUFF I64 (joint_0[0:0], i_0r1[0:0]);
  BUFF I65 (joint_0[1:1], i_0r1[1:1]);
  BUFF I66 (joint_0[2:2], i_0r1[2:2]);
  BUFF I67 (joint_0[3:3], i_0r1[3:3]);
  BUFF I68 (joint_0[4:4], i_0r1[4:4]);
  BUFF I69 (joint_0[5:5], i_0r1[5:5]);
  BUFF I70 (joint_0[6:6], i_0r1[6:6]);
  BUFF I71 (joint_0[7:7], i_0r1[7:7]);
  BUFF I72 (joint_0[8:8], i_0r1[8:8]);
  BUFF I73 (joint_0[9:9], i_0r1[9:9]);
  BUFF I74 (joint_0[10:10], i_0r1[10:10]);
  BUFF I75 (joint_0[11:11], i_0r1[11:11]);
  BUFF I76 (joint_0[12:12], i_0r1[12:12]);
  BUFF I77 (joint_0[13:13], i_0r1[13:13]);
  BUFF I78 (joint_0[14:14], i_0r1[14:14]);
  BUFF I79 (joint_0[15:15], i_0r1[15:15]);
  BUFF I80 (joint_0[16:16], i_0r1[16:16]);
  BUFF I81 (joint_0[17:17], i_0r1[17:17]);
  BUFF I82 (joint_0[18:18], i_0r1[18:18]);
  BUFF I83 (joint_0[19:19], i_0r1[19:19]);
  BUFF I84 (joint_0[20:20], i_0r1[20:20]);
  BUFF I85 (joint_0[21:21], i_0r1[21:21]);
  BUFF I86 (joint_0[22:22], i_0r1[22:22]);
  BUFF I87 (joint_0[23:23], i_0r1[23:23]);
  BUFF I88 (joint_0[24:24], i_0r1[24:24]);
  BUFF I89 (joint_0[25:25], i_0r1[25:25]);
  BUFF I90 (joint_0[26:26], i_0r1[26:26]);
  BUFF I91 (joint_0[27:27], i_0r1[27:27]);
  BUFF I92 (joint_0[28:28], i_0r1[28:28]);
  BUFF I93 (joint_0[29:29], i_0r1[29:29]);
  BUFF I94 (joint_0[30:30], i_0r1[30:30]);
  BUFF I95 (joint_0[31:31], i_0r1[31:31]);
  BUFF I96 (joint_0[32:32], i_1r1[0:0]);
  BUFF I97 (joint_0[33:33], i_1r1[1:1]);
  BUFF I98 (joint_0[34:34], i_1r1[2:2]);
  BUFF I99 (joint_0[35:35], i_1r1[3:3]);
  BUFF I100 (joint_0[36:36], i_1r1[4:4]);
  BUFF I101 (joint_0[37:37], i_1r1[5:5]);
  BUFF I102 (joint_0[38:38], i_1r1[6:6]);
  BUFF I103 (joint_0[39:39], i_1r1[7:7]);
  BUFF I104 (joint_0[40:40], i_1r1[8:8]);
  BUFF I105 (joint_0[41:41], i_1r1[9:9]);
  BUFF I106 (joint_0[42:42], i_1r1[10:10]);
  BUFF I107 (joint_0[43:43], i_1r1[11:11]);
  BUFF I108 (joint_0[44:44], i_1r1[12:12]);
  BUFF I109 (joint_0[45:45], i_1r1[13:13]);
  BUFF I110 (joint_0[46:46], i_1r1[14:14]);
  BUFF I111 (joint_0[47:47], i_1r1[15:15]);
  BUFF I112 (joint_0[48:48], i_1r1[16:16]);
  BUFF I113 (joint_0[49:49], i_1r1[17:17]);
  BUFF I114 (joint_0[50:50], i_1r1[18:18]);
  BUFF I115 (joint_0[51:51], i_1r1[19:19]);
  BUFF I116 (joint_0[52:52], i_1r1[20:20]);
  BUFF I117 (joint_0[53:53], i_1r1[21:21]);
  BUFF I118 (joint_0[54:54], i_1r1[22:22]);
  BUFF I119 (joint_0[55:55], i_1r1[23:23]);
  BUFF I120 (joint_0[56:56], i_1r1[24:24]);
  BUFF I121 (joint_0[57:57], i_1r1[25:25]);
  BUFF I122 (joint_0[58:58], i_1r1[26:26]);
  BUFF I123 (joint_0[59:59], i_1r1[27:27]);
  BUFF I124 (joint_0[60:60], i_1r1[28:28]);
  BUFF I125 (joint_0[61:61], i_1r1[29:29]);
  BUFF I126 (joint_0[62:62], i_1r1[30:30]);
  BUFF I127 (joint_0[63:63], i_1r1[31:31]);
  OR2 I128 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  C2 I129 (icomplete_0, i_2r, dcomplete_0);
  C2 I130 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I131 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I132 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I133 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I134 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I135 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I136 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I137 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I138 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I139 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I140 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I141 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I142 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I143 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I144 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I145 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I146 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I147 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I148 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I149 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I150 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I151 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I152 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I153 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I154 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I155 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I156 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I157 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I158 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I159 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I160 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I161 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I162 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I163 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I164 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I165 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I166 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I167 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I168 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I169 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I170 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I171 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I172 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I173 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I174 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I175 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I176 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I177 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I178 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I179 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I180 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I181 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I182 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I183 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I184 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I185 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I186 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I187 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I188 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I189 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I190 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I191 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I192 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I193 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I194 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I195 (o_0r1[1:1], joint_0[1:1]);
  BUFF I196 (o_0r1[2:2], joint_0[2:2]);
  BUFF I197 (o_0r1[3:3], joint_0[3:3]);
  BUFF I198 (o_0r1[4:4], joint_0[4:4]);
  BUFF I199 (o_0r1[5:5], joint_0[5:5]);
  BUFF I200 (o_0r1[6:6], joint_0[6:6]);
  BUFF I201 (o_0r1[7:7], joint_0[7:7]);
  BUFF I202 (o_0r1[8:8], joint_0[8:8]);
  BUFF I203 (o_0r1[9:9], joint_0[9:9]);
  BUFF I204 (o_0r1[10:10], joint_0[10:10]);
  BUFF I205 (o_0r1[11:11], joint_0[11:11]);
  BUFF I206 (o_0r1[12:12], joint_0[12:12]);
  BUFF I207 (o_0r1[13:13], joint_0[13:13]);
  BUFF I208 (o_0r1[14:14], joint_0[14:14]);
  BUFF I209 (o_0r1[15:15], joint_0[15:15]);
  BUFF I210 (o_0r1[16:16], joint_0[16:16]);
  BUFF I211 (o_0r1[17:17], joint_0[17:17]);
  BUFF I212 (o_0r1[18:18], joint_0[18:18]);
  BUFF I213 (o_0r1[19:19], joint_0[19:19]);
  BUFF I214 (o_0r1[20:20], joint_0[20:20]);
  BUFF I215 (o_0r1[21:21], joint_0[21:21]);
  BUFF I216 (o_0r1[22:22], joint_0[22:22]);
  BUFF I217 (o_0r1[23:23], joint_0[23:23]);
  BUFF I218 (o_0r1[24:24], joint_0[24:24]);
  BUFF I219 (o_0r1[25:25], joint_0[25:25]);
  BUFF I220 (o_0r1[26:26], joint_0[26:26]);
  BUFF I221 (o_0r1[27:27], joint_0[27:27]);
  BUFF I222 (o_0r1[28:28], joint_0[28:28]);
  BUFF I223 (o_0r1[29:29], joint_0[29:29]);
  BUFF I224 (o_0r1[30:30], joint_0[30:30]);
  BUFF I225 (o_0r1[31:31], joint_0[31:31]);
  BUFF I226 (o_0r1[32:32], joint_0[32:32]);
  BUFF I227 (o_0r1[33:33], joint_0[33:33]);
  BUFF I228 (o_0r1[34:34], joint_0[34:34]);
  BUFF I229 (o_0r1[35:35], joint_0[35:35]);
  BUFF I230 (o_0r1[36:36], joint_0[36:36]);
  BUFF I231 (o_0r1[37:37], joint_0[37:37]);
  BUFF I232 (o_0r1[38:38], joint_0[38:38]);
  BUFF I233 (o_0r1[39:39], joint_0[39:39]);
  BUFF I234 (o_0r1[40:40], joint_0[40:40]);
  BUFF I235 (o_0r1[41:41], joint_0[41:41]);
  BUFF I236 (o_0r1[42:42], joint_0[42:42]);
  BUFF I237 (o_0r1[43:43], joint_0[43:43]);
  BUFF I238 (o_0r1[44:44], joint_0[44:44]);
  BUFF I239 (o_0r1[45:45], joint_0[45:45]);
  BUFF I240 (o_0r1[46:46], joint_0[46:46]);
  BUFF I241 (o_0r1[47:47], joint_0[47:47]);
  BUFF I242 (o_0r1[48:48], joint_0[48:48]);
  BUFF I243 (o_0r1[49:49], joint_0[49:49]);
  BUFF I244 (o_0r1[50:50], joint_0[50:50]);
  BUFF I245 (o_0r1[51:51], joint_0[51:51]);
  BUFF I246 (o_0r1[52:52], joint_0[52:52]);
  BUFF I247 (o_0r1[53:53], joint_0[53:53]);
  BUFF I248 (o_0r1[54:54], joint_0[54:54]);
  BUFF I249 (o_0r1[55:55], joint_0[55:55]);
  BUFF I250 (o_0r1[56:56], joint_0[56:56]);
  BUFF I251 (o_0r1[57:57], joint_0[57:57]);
  BUFF I252 (o_0r1[58:58], joint_0[58:58]);
  BUFF I253 (o_0r1[59:59], joint_0[59:59]);
  BUFF I254 (o_0r1[60:60], joint_0[60:60]);
  BUFF I255 (o_0r1[61:61], joint_0[61:61]);
  BUFF I256 (o_0r1[62:62], joint_0[62:62]);
  BUFF I257 (o_0r1[63:63], joint_0[63:63]);
  BUFF I258 (i_0a, o_0a);
  BUFF I259 (i_1a, o_0a);
  BUFF I260 (i_2a, o_0a);
endmodule

// tko1m1_1nm1b1_2nei0w1bt1o0w1b TeakO [
//     (1,TeakOConstant 1 1),
//     (2,TeakOp TeakOpNotEqual [(0,0+:1),(1,0+:1)])] [One 1,One 1]
module tko1m1_1nm1b1_2nei0w1bt1o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire gocomp_0;
  wire termf_1;
  wire termt_1;
  wire xf2_0;
  wire xt2_0;
  wire [3:0] op2_0_0;
  OR2 I0 (gocomp_0, i_0r0, i_0r1);
  BUFF I1 (go_0, gocomp_0);
  BUFF I2 (termt_1, go_0);
  GND I3 (termf_1);
  C2 I4 (op2_0_0[0:0], termf_1, i_0r0);
  C2 I5 (op2_0_0[1:1], termf_1, i_0r1);
  C2 I6 (op2_0_0[2:2], termt_1, i_0r0);
  C2 I7 (op2_0_0[3:3], termt_1, i_0r1);
  OR2 I8 (xf2_0, op2_0_0[1:1], op2_0_0[2:2]);
  OR2 I9 (xt2_0, op2_0_0[0:0], op2_0_0[3:3]);
  BUFF I10 (o_0r1, xf2_0);
  BUFF I11 (o_0r0, xt2_0);
  BUFF I12 (i_0a, o_0a);
endmodule

// tko1m1_1nm1b1_2eqi0w1bt1o0w1b TeakO [
//     (1,TeakOConstant 1 1),
//     (2,TeakOp TeakOpEqual [(0,0+:1),(1,0+:1)])] [One 1,One 1]
module tko1m1_1nm1b1_2eqi0w1bt1o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire gocomp_0;
  wire termf_1;
  wire termt_1;
  wire xf2_0;
  wire xt2_0;
  wire [3:0] op2_0_0;
  OR2 I0 (gocomp_0, i_0r0, i_0r1);
  BUFF I1 (go_0, gocomp_0);
  BUFF I2 (termt_1, go_0);
  GND I3 (termf_1);
  C2 I4 (op2_0_0[0:0], termf_1, i_0r0);
  C2 I5 (op2_0_0[1:1], termf_1, i_0r1);
  C2 I6 (op2_0_0[2:2], termt_1, i_0r0);
  C2 I7 (op2_0_0[3:3], termt_1, i_0r1);
  OR2 I8 (xf2_0, op2_0_0[1:1], op2_0_0[2:2]);
  OR2 I9 (xt2_0, op2_0_0[0:0], op2_0_0[3:3]);
  BUFF I10 (o_0r0, xf2_0);
  BUFF I11 (o_0r1, xt2_0);
  BUFF I12 (i_0a, o_0a);
endmodule

// tko3m4_1nm1b0_2api0w3bt1o0w1b_3nm4b1_4addt2o0w4bt3o0w4b TeakO [
//     (1,TeakOConstant 1 0),
//     (2,TeakOAppend 1 [(0,0+:3),(1,0+:1)]),
//     (3,TeakOConstant 4 1),
//     (4,TeakOp TeakOpAdd [(2,0+:4),(3,0+:4)])] [One 3,One 4]
module tko3m4_1nm1b0_2api0w3bt1o0w1b_3nm4b1_4addt2o0w4bt3o0w4b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [2:0] gocomp_0;
  wire termf_1;
  wire [3:0] termf_2;
  wire [3:0] termf_3;
  wire termt_1;
  wire [3:0] termt_2;
  wire [3:0] termt_3;
  wire [3:0] cf4__0;
  wire [3:0] ct4__0;
  wire [3:0] ha4__0;
  wire [7:0] fa4_1min_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [7:0] fa4_2min_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [7:0] fa4_3min_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I3 (go_0, gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  BUFF I4 (termf_1, go_0);
  GND I5 (termt_1);
  BUFF I6 (termf_2[0:0], i_0r0[0:0]);
  BUFF I7 (termf_2[1:1], i_0r0[1:1]);
  BUFF I8 (termf_2[2:2], i_0r0[2:2]);
  BUFF I9 (termf_2[3:3], termf_1);
  BUFF I10 (termt_2[0:0], i_0r1[0:0]);
  BUFF I11 (termt_2[1:1], i_0r1[1:1]);
  BUFF I12 (termt_2[2:2], i_0r1[2:2]);
  BUFF I13 (termt_2[3:3], termt_1);
  BUFF I14 (termt_3[0:0], go_0);
  GND I15 (termf_3[0:0]);
  BUFF I16 (termf_3[1:1], go_0);
  BUFF I17 (termf_3[2:2], go_0);
  BUFF I18 (termf_3[3:3], go_0);
  GND I19 (termt_3[1:1]);
  GND I20 (termt_3[2:2]);
  GND I21 (termt_3[3:3]);
  C2 I22 (ha4__0[0:0], termf_3[0:0], termf_2[0:0]);
  C2 I23 (ha4__0[1:1], termf_3[0:0], termt_2[0:0]);
  C2 I24 (ha4__0[2:2], termt_3[0:0], termf_2[0:0]);
  C2 I25 (ha4__0[3:3], termt_3[0:0], termt_2[0:0]);
  OR3 I26 (cf4__0[0:0], ha4__0[0:0], ha4__0[1:1], ha4__0[2:2]);
  BUFF I27 (ct4__0[0:0], ha4__0[3:3]);
  OR2 I28 (o_0r0[0:0], ha4__0[0:0], ha4__0[3:3]);
  OR2 I29 (o_0r1[0:0], ha4__0[1:1], ha4__0[2:2]);
  C3 I30 (fa4_1min_0[0:0], cf4__0[0:0], termf_3[1:1], termf_2[1:1]);
  C3 I31 (fa4_1min_0[1:1], cf4__0[0:0], termf_3[1:1], termt_2[1:1]);
  C3 I32 (fa4_1min_0[2:2], cf4__0[0:0], termt_3[1:1], termf_2[1:1]);
  C3 I33 (fa4_1min_0[3:3], cf4__0[0:0], termt_3[1:1], termt_2[1:1]);
  C3 I34 (fa4_1min_0[4:4], ct4__0[0:0], termf_3[1:1], termf_2[1:1]);
  C3 I35 (fa4_1min_0[5:5], ct4__0[0:0], termf_3[1:1], termt_2[1:1]);
  C3 I36 (fa4_1min_0[6:6], ct4__0[0:0], termt_3[1:1], termf_2[1:1]);
  C3 I37 (fa4_1min_0[7:7], ct4__0[0:0], termt_3[1:1], termt_2[1:1]);
  NOR3 I38 (simp471_0[0:0], fa4_1min_0[0:0], fa4_1min_0[3:3], fa4_1min_0[5:5]);
  INV I39 (simp471_0[1:1], fa4_1min_0[6:6]);
  NAND2 I40 (o_0r0[1:1], simp471_0[0:0], simp471_0[1:1]);
  NOR3 I41 (simp481_0[0:0], fa4_1min_0[1:1], fa4_1min_0[2:2], fa4_1min_0[4:4]);
  INV I42 (simp481_0[1:1], fa4_1min_0[7:7]);
  NAND2 I43 (o_0r1[1:1], simp481_0[0:0], simp481_0[1:1]);
  AO222 I44 (ct4__0[1:1], termt_2[1:1], termt_3[1:1], termt_2[1:1], ct4__0[0:0], termt_3[1:1], ct4__0[0:0]);
  AO222 I45 (cf4__0[1:1], termf_2[1:1], termf_3[1:1], termf_2[1:1], cf4__0[0:0], termf_3[1:1], cf4__0[0:0]);
  C3 I46 (fa4_2min_0[0:0], cf4__0[1:1], termf_3[2:2], termf_2[2:2]);
  C3 I47 (fa4_2min_0[1:1], cf4__0[1:1], termf_3[2:2], termt_2[2:2]);
  C3 I48 (fa4_2min_0[2:2], cf4__0[1:1], termt_3[2:2], termf_2[2:2]);
  C3 I49 (fa4_2min_0[3:3], cf4__0[1:1], termt_3[2:2], termt_2[2:2]);
  C3 I50 (fa4_2min_0[4:4], ct4__0[1:1], termf_3[2:2], termf_2[2:2]);
  C3 I51 (fa4_2min_0[5:5], ct4__0[1:1], termf_3[2:2], termt_2[2:2]);
  C3 I52 (fa4_2min_0[6:6], ct4__0[1:1], termt_3[2:2], termf_2[2:2]);
  C3 I53 (fa4_2min_0[7:7], ct4__0[1:1], termt_3[2:2], termt_2[2:2]);
  NOR3 I54 (simp601_0[0:0], fa4_2min_0[0:0], fa4_2min_0[3:3], fa4_2min_0[5:5]);
  INV I55 (simp601_0[1:1], fa4_2min_0[6:6]);
  NAND2 I56 (o_0r0[2:2], simp601_0[0:0], simp601_0[1:1]);
  NOR3 I57 (simp611_0[0:0], fa4_2min_0[1:1], fa4_2min_0[2:2], fa4_2min_0[4:4]);
  INV I58 (simp611_0[1:1], fa4_2min_0[7:7]);
  NAND2 I59 (o_0r1[2:2], simp611_0[0:0], simp611_0[1:1]);
  AO222 I60 (ct4__0[2:2], termt_2[2:2], termt_3[2:2], termt_2[2:2], ct4__0[1:1], termt_3[2:2], ct4__0[1:1]);
  AO222 I61 (cf4__0[2:2], termf_2[2:2], termf_3[2:2], termf_2[2:2], cf4__0[1:1], termf_3[2:2], cf4__0[1:1]);
  C3 I62 (fa4_3min_0[0:0], cf4__0[2:2], termf_3[3:3], termf_2[3:3]);
  C3 I63 (fa4_3min_0[1:1], cf4__0[2:2], termf_3[3:3], termt_2[3:3]);
  C3 I64 (fa4_3min_0[2:2], cf4__0[2:2], termt_3[3:3], termf_2[3:3]);
  C3 I65 (fa4_3min_0[3:3], cf4__0[2:2], termt_3[3:3], termt_2[3:3]);
  C3 I66 (fa4_3min_0[4:4], ct4__0[2:2], termf_3[3:3], termf_2[3:3]);
  C3 I67 (fa4_3min_0[5:5], ct4__0[2:2], termf_3[3:3], termt_2[3:3]);
  C3 I68 (fa4_3min_0[6:6], ct4__0[2:2], termt_3[3:3], termf_2[3:3]);
  C3 I69 (fa4_3min_0[7:7], ct4__0[2:2], termt_3[3:3], termt_2[3:3]);
  NOR3 I70 (simp731_0[0:0], fa4_3min_0[0:0], fa4_3min_0[3:3], fa4_3min_0[5:5]);
  INV I71 (simp731_0[1:1], fa4_3min_0[6:6]);
  NAND2 I72 (o_0r0[3:3], simp731_0[0:0], simp731_0[1:1]);
  NOR3 I73 (simp741_0[0:0], fa4_3min_0[1:1], fa4_3min_0[2:2], fa4_3min_0[4:4]);
  INV I74 (simp741_0[1:1], fa4_3min_0[7:7]);
  NAND2 I75 (o_0r1[3:3], simp741_0[0:0], simp741_0[1:1]);
  AO222 I76 (ct4__0[3:3], termt_2[3:3], termt_3[3:3], termt_2[3:3], ct4__0[2:2], termt_3[3:3], ct4__0[2:2]);
  AO222 I77 (cf4__0[3:3], termf_2[3:3], termf_3[3:3], termf_2[3:3], cf4__0[2:2], termf_3[3:3], cf4__0[2:2]);
  BUFF I78 (i_0a, o_0a);
endmodule

// tko32m1_1nm32b0_2sgti0w32bt1o0w32b TeakO [
//     (1,TeakOConstant 32 0),
//     (2,TeakOp TeakOpSignedGT [(0,0+:32),(1,0+:32)])] [One 32,One 1]
module tko32m1_1nm32b0_2sgti0w32bt1o0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [31:0] gocomp_0;
  wire [10:0] simp341_0;
  wire [3:0] simp342_0;
  wire [1:0] simp343_0;
  wire [31:0] termf_1;
  wire [31:0] termt_1;
  wire [31:0] eq2_0;
  wire [31:0] gt2_0;
  wire [31:0] lt2_0;
  wire oeq2_0;
  wire ogt2_0;
  wire olt2_0;
  wire [31:0] mt0_2_0;
  wire [31:0] mt3_2_0;
  wire [15:0] comb2o_0;
  wire [15:0] comb2o_1;
  wire [15:0] comb2o_2;
  wire [7:0] comb2ro_0;
  wire [7:0] comb2ro_1;
  wire [7:0] comb2ro_2;
  wire [3:0] comb2rro_0;
  wire [3:0] comb2rro_1;
  wire [3:0] comb2rro_2;
  wire [1:0] comb2rrro_0;
  wire [1:0] comb2rrro_1;
  wire [1:0] comb2rrro_2;
  wire comb2rrrr0ltint_0;
  wire comb2rrrr0gtint_0;
  wire comb2rrr0ltint_0;
  wire comb2rrr0gtint_0;
  wire comb2rrr1ltint_0;
  wire comb2rrr1gtint_0;
  wire comb2rr0ltint_0;
  wire comb2rr0gtint_0;
  wire comb2rr1ltint_0;
  wire comb2rr1gtint_0;
  wire comb2rr2ltint_0;
  wire comb2rr2gtint_0;
  wire comb2rr3ltint_0;
  wire comb2rr3gtint_0;
  wire comb2r0ltint_0;
  wire comb2r0gtint_0;
  wire comb2r1ltint_0;
  wire comb2r1gtint_0;
  wire comb2r2ltint_0;
  wire comb2r2gtint_0;
  wire comb2r3ltint_0;
  wire comb2r3gtint_0;
  wire comb2r4ltint_0;
  wire comb2r4gtint_0;
  wire comb2r5ltint_0;
  wire comb2r5gtint_0;
  wire comb2r6ltint_0;
  wire comb2r6gtint_0;
  wire comb2r7ltint_0;
  wire comb2r7gtint_0;
  wire comb20ltint_0;
  wire comb20gtint_0;
  wire comb21ltint_0;
  wire comb21gtint_0;
  wire comb22ltint_0;
  wire comb22gtint_0;
  wire comb23ltint_0;
  wire comb23gtint_0;
  wire comb24ltint_0;
  wire comb24gtint_0;
  wire comb25ltint_0;
  wire comb25gtint_0;
  wire comb26ltint_0;
  wire comb26gtint_0;
  wire comb27ltint_0;
  wire comb27gtint_0;
  wire comb28ltint_0;
  wire comb28gtint_0;
  wire comb29ltint_0;
  wire comb29gtint_0;
  wire comb210ltint_0;
  wire comb210gtint_0;
  wire comb211ltint_0;
  wire comb211gtint_0;
  wire comb212ltint_0;
  wire comb212gtint_0;
  wire comb213ltint_0;
  wire comb213gtint_0;
  wire comb214ltint_0;
  wire comb214gtint_0;
  wire comb215ltint_0;
  wire comb215gtint_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I32 (simp341_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I33 (simp341_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I34 (simp341_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I35 (simp341_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I36 (simp341_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I37 (simp341_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I38 (simp341_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I39 (simp341_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I40 (simp341_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I41 (simp341_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C2 I42 (simp341_0[10:10], gocomp_0[30:30], gocomp_0[31:31]);
  C3 I43 (simp342_0[0:0], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  C3 I44 (simp342_0[1:1], simp341_0[3:3], simp341_0[4:4], simp341_0[5:5]);
  C3 I45 (simp342_0[2:2], simp341_0[6:6], simp341_0[7:7], simp341_0[8:8]);
  C2 I46 (simp342_0[3:3], simp341_0[9:9], simp341_0[10:10]);
  C3 I47 (simp343_0[0:0], simp342_0[0:0], simp342_0[1:1], simp342_0[2:2]);
  BUFF I48 (simp343_0[1:1], simp342_0[3:3]);
  C2 I49 (go_0, simp343_0[0:0], simp343_0[1:1]);
  BUFF I50 (termf_1[0:0], go_0);
  BUFF I51 (termf_1[1:1], go_0);
  BUFF I52 (termf_1[2:2], go_0);
  BUFF I53 (termf_1[3:3], go_0);
  BUFF I54 (termf_1[4:4], go_0);
  BUFF I55 (termf_1[5:5], go_0);
  BUFF I56 (termf_1[6:6], go_0);
  BUFF I57 (termf_1[7:7], go_0);
  BUFF I58 (termf_1[8:8], go_0);
  BUFF I59 (termf_1[9:9], go_0);
  BUFF I60 (termf_1[10:10], go_0);
  BUFF I61 (termf_1[11:11], go_0);
  BUFF I62 (termf_1[12:12], go_0);
  BUFF I63 (termf_1[13:13], go_0);
  BUFF I64 (termf_1[14:14], go_0);
  BUFF I65 (termf_1[15:15], go_0);
  BUFF I66 (termf_1[16:16], go_0);
  BUFF I67 (termf_1[17:17], go_0);
  BUFF I68 (termf_1[18:18], go_0);
  BUFF I69 (termf_1[19:19], go_0);
  BUFF I70 (termf_1[20:20], go_0);
  BUFF I71 (termf_1[21:21], go_0);
  BUFF I72 (termf_1[22:22], go_0);
  BUFF I73 (termf_1[23:23], go_0);
  BUFF I74 (termf_1[24:24], go_0);
  BUFF I75 (termf_1[25:25], go_0);
  BUFF I76 (termf_1[26:26], go_0);
  BUFF I77 (termf_1[27:27], go_0);
  BUFF I78 (termf_1[28:28], go_0);
  BUFF I79 (termf_1[29:29], go_0);
  BUFF I80 (termf_1[30:30], go_0);
  BUFF I81 (termf_1[31:31], go_0);
  GND I82 (termt_1[0:0]);
  GND I83 (termt_1[1:1]);
  GND I84 (termt_1[2:2]);
  GND I85 (termt_1[3:3]);
  GND I86 (termt_1[4:4]);
  GND I87 (termt_1[5:5]);
  GND I88 (termt_1[6:6]);
  GND I89 (termt_1[7:7]);
  GND I90 (termt_1[8:8]);
  GND I91 (termt_1[9:9]);
  GND I92 (termt_1[10:10]);
  GND I93 (termt_1[11:11]);
  GND I94 (termt_1[12:12]);
  GND I95 (termt_1[13:13]);
  GND I96 (termt_1[14:14]);
  GND I97 (termt_1[15:15]);
  GND I98 (termt_1[16:16]);
  GND I99 (termt_1[17:17]);
  GND I100 (termt_1[18:18]);
  GND I101 (termt_1[19:19]);
  GND I102 (termt_1[20:20]);
  GND I103 (termt_1[21:21]);
  GND I104 (termt_1[22:22]);
  GND I105 (termt_1[23:23]);
  GND I106 (termt_1[24:24]);
  GND I107 (termt_1[25:25]);
  GND I108 (termt_1[26:26]);
  GND I109 (termt_1[27:27]);
  GND I110 (termt_1[28:28]);
  GND I111 (termt_1[29:29]);
  GND I112 (termt_1[30:30]);
  GND I113 (termt_1[31:31]);
  C2 I114 (mt0_2_0[0:0], i_0r0[0:0], termf_1[0:0]);
  C2 I115 (mt0_2_0[1:1], i_0r0[1:1], termf_1[1:1]);
  C2 I116 (mt0_2_0[2:2], i_0r0[2:2], termf_1[2:2]);
  C2 I117 (mt0_2_0[3:3], i_0r0[3:3], termf_1[3:3]);
  C2 I118 (mt0_2_0[4:4], i_0r0[4:4], termf_1[4:4]);
  C2 I119 (mt0_2_0[5:5], i_0r0[5:5], termf_1[5:5]);
  C2 I120 (mt0_2_0[6:6], i_0r0[6:6], termf_1[6:6]);
  C2 I121 (mt0_2_0[7:7], i_0r0[7:7], termf_1[7:7]);
  C2 I122 (mt0_2_0[8:8], i_0r0[8:8], termf_1[8:8]);
  C2 I123 (mt0_2_0[9:9], i_0r0[9:9], termf_1[9:9]);
  C2 I124 (mt0_2_0[10:10], i_0r0[10:10], termf_1[10:10]);
  C2 I125 (mt0_2_0[11:11], i_0r0[11:11], termf_1[11:11]);
  C2 I126 (mt0_2_0[12:12], i_0r0[12:12], termf_1[12:12]);
  C2 I127 (mt0_2_0[13:13], i_0r0[13:13], termf_1[13:13]);
  C2 I128 (mt0_2_0[14:14], i_0r0[14:14], termf_1[14:14]);
  C2 I129 (mt0_2_0[15:15], i_0r0[15:15], termf_1[15:15]);
  C2 I130 (mt0_2_0[16:16], i_0r0[16:16], termf_1[16:16]);
  C2 I131 (mt0_2_0[17:17], i_0r0[17:17], termf_1[17:17]);
  C2 I132 (mt0_2_0[18:18], i_0r0[18:18], termf_1[18:18]);
  C2 I133 (mt0_2_0[19:19], i_0r0[19:19], termf_1[19:19]);
  C2 I134 (mt0_2_0[20:20], i_0r0[20:20], termf_1[20:20]);
  C2 I135 (mt0_2_0[21:21], i_0r0[21:21], termf_1[21:21]);
  C2 I136 (mt0_2_0[22:22], i_0r0[22:22], termf_1[22:22]);
  C2 I137 (mt0_2_0[23:23], i_0r0[23:23], termf_1[23:23]);
  C2 I138 (mt0_2_0[24:24], i_0r0[24:24], termf_1[24:24]);
  C2 I139 (mt0_2_0[25:25], i_0r0[25:25], termf_1[25:25]);
  C2 I140 (mt0_2_0[26:26], i_0r0[26:26], termf_1[26:26]);
  C2 I141 (mt0_2_0[27:27], i_0r0[27:27], termf_1[27:27]);
  C2 I142 (mt0_2_0[28:28], i_0r0[28:28], termf_1[28:28]);
  C2 I143 (mt0_2_0[29:29], i_0r0[29:29], termf_1[29:29]);
  C2 I144 (mt0_2_0[30:30], i_0r0[30:30], termf_1[30:30]);
  C2 I145 (mt0_2_0[31:31], i_0r0[31:31], termf_1[31:31]);
  C2 I146 (mt3_2_0[0:0], i_0r1[0:0], termt_1[0:0]);
  C2 I147 (mt3_2_0[1:1], i_0r1[1:1], termt_1[1:1]);
  C2 I148 (mt3_2_0[2:2], i_0r1[2:2], termt_1[2:2]);
  C2 I149 (mt3_2_0[3:3], i_0r1[3:3], termt_1[3:3]);
  C2 I150 (mt3_2_0[4:4], i_0r1[4:4], termt_1[4:4]);
  C2 I151 (mt3_2_0[5:5], i_0r1[5:5], termt_1[5:5]);
  C2 I152 (mt3_2_0[6:6], i_0r1[6:6], termt_1[6:6]);
  C2 I153 (mt3_2_0[7:7], i_0r1[7:7], termt_1[7:7]);
  C2 I154 (mt3_2_0[8:8], i_0r1[8:8], termt_1[8:8]);
  C2 I155 (mt3_2_0[9:9], i_0r1[9:9], termt_1[9:9]);
  C2 I156 (mt3_2_0[10:10], i_0r1[10:10], termt_1[10:10]);
  C2 I157 (mt3_2_0[11:11], i_0r1[11:11], termt_1[11:11]);
  C2 I158 (mt3_2_0[12:12], i_0r1[12:12], termt_1[12:12]);
  C2 I159 (mt3_2_0[13:13], i_0r1[13:13], termt_1[13:13]);
  C2 I160 (mt3_2_0[14:14], i_0r1[14:14], termt_1[14:14]);
  C2 I161 (mt3_2_0[15:15], i_0r1[15:15], termt_1[15:15]);
  C2 I162 (mt3_2_0[16:16], i_0r1[16:16], termt_1[16:16]);
  C2 I163 (mt3_2_0[17:17], i_0r1[17:17], termt_1[17:17]);
  C2 I164 (mt3_2_0[18:18], i_0r1[18:18], termt_1[18:18]);
  C2 I165 (mt3_2_0[19:19], i_0r1[19:19], termt_1[19:19]);
  C2 I166 (mt3_2_0[20:20], i_0r1[20:20], termt_1[20:20]);
  C2 I167 (mt3_2_0[21:21], i_0r1[21:21], termt_1[21:21]);
  C2 I168 (mt3_2_0[22:22], i_0r1[22:22], termt_1[22:22]);
  C2 I169 (mt3_2_0[23:23], i_0r1[23:23], termt_1[23:23]);
  C2 I170 (mt3_2_0[24:24], i_0r1[24:24], termt_1[24:24]);
  C2 I171 (mt3_2_0[25:25], i_0r1[25:25], termt_1[25:25]);
  C2 I172 (mt3_2_0[26:26], i_0r1[26:26], termt_1[26:26]);
  C2 I173 (mt3_2_0[27:27], i_0r1[27:27], termt_1[27:27]);
  C2 I174 (mt3_2_0[28:28], i_0r1[28:28], termt_1[28:28]);
  C2 I175 (mt3_2_0[29:29], i_0r1[29:29], termt_1[29:29]);
  C2 I176 (mt3_2_0[30:30], i_0r1[30:30], termt_1[30:30]);
  C2 I177 (mt3_2_0[31:31], i_0r1[31:31], termt_1[31:31]);
  C2 I178 (lt2_0[0:0], i_0r0[0:0], termt_1[0:0]);
  C2 I179 (lt2_0[1:1], i_0r0[1:1], termt_1[1:1]);
  C2 I180 (lt2_0[2:2], i_0r0[2:2], termt_1[2:2]);
  C2 I181 (lt2_0[3:3], i_0r0[3:3], termt_1[3:3]);
  C2 I182 (lt2_0[4:4], i_0r0[4:4], termt_1[4:4]);
  C2 I183 (lt2_0[5:5], i_0r0[5:5], termt_1[5:5]);
  C2 I184 (lt2_0[6:6], i_0r0[6:6], termt_1[6:6]);
  C2 I185 (lt2_0[7:7], i_0r0[7:7], termt_1[7:7]);
  C2 I186 (lt2_0[8:8], i_0r0[8:8], termt_1[8:8]);
  C2 I187 (lt2_0[9:9], i_0r0[9:9], termt_1[9:9]);
  C2 I188 (lt2_0[10:10], i_0r0[10:10], termt_1[10:10]);
  C2 I189 (lt2_0[11:11], i_0r0[11:11], termt_1[11:11]);
  C2 I190 (lt2_0[12:12], i_0r0[12:12], termt_1[12:12]);
  C2 I191 (lt2_0[13:13], i_0r0[13:13], termt_1[13:13]);
  C2 I192 (lt2_0[14:14], i_0r0[14:14], termt_1[14:14]);
  C2 I193 (lt2_0[15:15], i_0r0[15:15], termt_1[15:15]);
  C2 I194 (lt2_0[16:16], i_0r0[16:16], termt_1[16:16]);
  C2 I195 (lt2_0[17:17], i_0r0[17:17], termt_1[17:17]);
  C2 I196 (lt2_0[18:18], i_0r0[18:18], termt_1[18:18]);
  C2 I197 (lt2_0[19:19], i_0r0[19:19], termt_1[19:19]);
  C2 I198 (lt2_0[20:20], i_0r0[20:20], termt_1[20:20]);
  C2 I199 (lt2_0[21:21], i_0r0[21:21], termt_1[21:21]);
  C2 I200 (lt2_0[22:22], i_0r0[22:22], termt_1[22:22]);
  C2 I201 (lt2_0[23:23], i_0r0[23:23], termt_1[23:23]);
  C2 I202 (lt2_0[24:24], i_0r0[24:24], termt_1[24:24]);
  C2 I203 (lt2_0[25:25], i_0r0[25:25], termt_1[25:25]);
  C2 I204 (lt2_0[26:26], i_0r0[26:26], termt_1[26:26]);
  C2 I205 (lt2_0[27:27], i_0r0[27:27], termt_1[27:27]);
  C2 I206 (lt2_0[28:28], i_0r0[28:28], termt_1[28:28]);
  C2 I207 (lt2_0[29:29], i_0r0[29:29], termt_1[29:29]);
  C2 I208 (lt2_0[30:30], i_0r0[30:30], termt_1[30:30]);
  C2 I209 (lt2_0[31:31], i_0r0[31:31], termt_1[31:31]);
  C2 I210 (gt2_0[0:0], i_0r1[0:0], termf_1[0:0]);
  C2 I211 (gt2_0[1:1], i_0r1[1:1], termf_1[1:1]);
  C2 I212 (gt2_0[2:2], i_0r1[2:2], termf_1[2:2]);
  C2 I213 (gt2_0[3:3], i_0r1[3:3], termf_1[3:3]);
  C2 I214 (gt2_0[4:4], i_0r1[4:4], termf_1[4:4]);
  C2 I215 (gt2_0[5:5], i_0r1[5:5], termf_1[5:5]);
  C2 I216 (gt2_0[6:6], i_0r1[6:6], termf_1[6:6]);
  C2 I217 (gt2_0[7:7], i_0r1[7:7], termf_1[7:7]);
  C2 I218 (gt2_0[8:8], i_0r1[8:8], termf_1[8:8]);
  C2 I219 (gt2_0[9:9], i_0r1[9:9], termf_1[9:9]);
  C2 I220 (gt2_0[10:10], i_0r1[10:10], termf_1[10:10]);
  C2 I221 (gt2_0[11:11], i_0r1[11:11], termf_1[11:11]);
  C2 I222 (gt2_0[12:12], i_0r1[12:12], termf_1[12:12]);
  C2 I223 (gt2_0[13:13], i_0r1[13:13], termf_1[13:13]);
  C2 I224 (gt2_0[14:14], i_0r1[14:14], termf_1[14:14]);
  C2 I225 (gt2_0[15:15], i_0r1[15:15], termf_1[15:15]);
  C2 I226 (gt2_0[16:16], i_0r1[16:16], termf_1[16:16]);
  C2 I227 (gt2_0[17:17], i_0r1[17:17], termf_1[17:17]);
  C2 I228 (gt2_0[18:18], i_0r1[18:18], termf_1[18:18]);
  C2 I229 (gt2_0[19:19], i_0r1[19:19], termf_1[19:19]);
  C2 I230 (gt2_0[20:20], i_0r1[20:20], termf_1[20:20]);
  C2 I231 (gt2_0[21:21], i_0r1[21:21], termf_1[21:21]);
  C2 I232 (gt2_0[22:22], i_0r1[22:22], termf_1[22:22]);
  C2 I233 (gt2_0[23:23], i_0r1[23:23], termf_1[23:23]);
  C2 I234 (gt2_0[24:24], i_0r1[24:24], termf_1[24:24]);
  C2 I235 (gt2_0[25:25], i_0r1[25:25], termf_1[25:25]);
  C2 I236 (gt2_0[26:26], i_0r1[26:26], termf_1[26:26]);
  C2 I237 (gt2_0[27:27], i_0r1[27:27], termf_1[27:27]);
  C2 I238 (gt2_0[28:28], i_0r1[28:28], termf_1[28:28]);
  C2 I239 (gt2_0[29:29], i_0r1[29:29], termf_1[29:29]);
  C2 I240 (gt2_0[30:30], i_0r1[30:30], termf_1[30:30]);
  C2 I241 (gt2_0[31:31], i_0r1[31:31], termf_1[31:31]);
  OR2 I242 (eq2_0[0:0], mt0_2_0[0:0], mt3_2_0[0:0]);
  OR2 I243 (eq2_0[1:1], mt0_2_0[1:1], mt3_2_0[1:1]);
  OR2 I244 (eq2_0[2:2], mt0_2_0[2:2], mt3_2_0[2:2]);
  OR2 I245 (eq2_0[3:3], mt0_2_0[3:3], mt3_2_0[3:3]);
  OR2 I246 (eq2_0[4:4], mt0_2_0[4:4], mt3_2_0[4:4]);
  OR2 I247 (eq2_0[5:5], mt0_2_0[5:5], mt3_2_0[5:5]);
  OR2 I248 (eq2_0[6:6], mt0_2_0[6:6], mt3_2_0[6:6]);
  OR2 I249 (eq2_0[7:7], mt0_2_0[7:7], mt3_2_0[7:7]);
  OR2 I250 (eq2_0[8:8], mt0_2_0[8:8], mt3_2_0[8:8]);
  OR2 I251 (eq2_0[9:9], mt0_2_0[9:9], mt3_2_0[9:9]);
  OR2 I252 (eq2_0[10:10], mt0_2_0[10:10], mt3_2_0[10:10]);
  OR2 I253 (eq2_0[11:11], mt0_2_0[11:11], mt3_2_0[11:11]);
  OR2 I254 (eq2_0[12:12], mt0_2_0[12:12], mt3_2_0[12:12]);
  OR2 I255 (eq2_0[13:13], mt0_2_0[13:13], mt3_2_0[13:13]);
  OR2 I256 (eq2_0[14:14], mt0_2_0[14:14], mt3_2_0[14:14]);
  OR2 I257 (eq2_0[15:15], mt0_2_0[15:15], mt3_2_0[15:15]);
  OR2 I258 (eq2_0[16:16], mt0_2_0[16:16], mt3_2_0[16:16]);
  OR2 I259 (eq2_0[17:17], mt0_2_0[17:17], mt3_2_0[17:17]);
  OR2 I260 (eq2_0[18:18], mt0_2_0[18:18], mt3_2_0[18:18]);
  OR2 I261 (eq2_0[19:19], mt0_2_0[19:19], mt3_2_0[19:19]);
  OR2 I262 (eq2_0[20:20], mt0_2_0[20:20], mt3_2_0[20:20]);
  OR2 I263 (eq2_0[21:21], mt0_2_0[21:21], mt3_2_0[21:21]);
  OR2 I264 (eq2_0[22:22], mt0_2_0[22:22], mt3_2_0[22:22]);
  OR2 I265 (eq2_0[23:23], mt0_2_0[23:23], mt3_2_0[23:23]);
  OR2 I266 (eq2_0[24:24], mt0_2_0[24:24], mt3_2_0[24:24]);
  OR2 I267 (eq2_0[25:25], mt0_2_0[25:25], mt3_2_0[25:25]);
  OR2 I268 (eq2_0[26:26], mt0_2_0[26:26], mt3_2_0[26:26]);
  OR2 I269 (eq2_0[27:27], mt0_2_0[27:27], mt3_2_0[27:27]);
  OR2 I270 (eq2_0[28:28], mt0_2_0[28:28], mt3_2_0[28:28]);
  OR2 I271 (eq2_0[29:29], mt0_2_0[29:29], mt3_2_0[29:29]);
  OR2 I272 (eq2_0[30:30], mt0_2_0[30:30], mt3_2_0[30:30]);
  OR2 I273 (eq2_0[31:31], mt0_2_0[31:31], mt3_2_0[31:31]);
  C2 I274 (oeq2_0, comb2rrro_0[0:0], comb2rrro_0[1:1]);
  C2 I275 (comb2rrrr0ltint_0, comb2rrro_1[0:0], comb2rrro_0[1:1]);
  C2 I276 (comb2rrrr0gtint_0, comb2rrro_2[0:0], comb2rrro_0[1:1]);
  OR2 I277 (olt2_0, comb2rrrr0ltint_0, comb2rrro_1[1:1]);
  OR2 I278 (ogt2_0, comb2rrrr0gtint_0, comb2rrro_2[1:1]);
  C2 I279 (comb2rrro_0[0:0], comb2rro_0[0:0], comb2rro_0[1:1]);
  C2 I280 (comb2rrr0ltint_0, comb2rro_1[0:0], comb2rro_0[1:1]);
  C2 I281 (comb2rrr0gtint_0, comb2rro_2[0:0], comb2rro_0[1:1]);
  OR2 I282 (comb2rrro_1[0:0], comb2rrr0ltint_0, comb2rro_1[1:1]);
  OR2 I283 (comb2rrro_2[0:0], comb2rrr0gtint_0, comb2rro_2[1:1]);
  C2 I284 (comb2rrro_0[1:1], comb2rro_0[2:2], comb2rro_0[3:3]);
  C2 I285 (comb2rrr1ltint_0, comb2rro_1[2:2], comb2rro_0[3:3]);
  C2 I286 (comb2rrr1gtint_0, comb2rro_2[2:2], comb2rro_0[3:3]);
  OR2 I287 (comb2rrro_1[1:1], comb2rrr1ltint_0, comb2rro_1[3:3]);
  OR2 I288 (comb2rrro_2[1:1], comb2rrr1gtint_0, comb2rro_2[3:3]);
  C2 I289 (comb2rro_0[0:0], comb2ro_0[0:0], comb2ro_0[1:1]);
  C2 I290 (comb2rr0ltint_0, comb2ro_1[0:0], comb2ro_0[1:1]);
  C2 I291 (comb2rr0gtint_0, comb2ro_2[0:0], comb2ro_0[1:1]);
  OR2 I292 (comb2rro_1[0:0], comb2rr0ltint_0, comb2ro_1[1:1]);
  OR2 I293 (comb2rro_2[0:0], comb2rr0gtint_0, comb2ro_2[1:1]);
  C2 I294 (comb2rro_0[1:1], comb2ro_0[2:2], comb2ro_0[3:3]);
  C2 I295 (comb2rr1ltint_0, comb2ro_1[2:2], comb2ro_0[3:3]);
  C2 I296 (comb2rr1gtint_0, comb2ro_2[2:2], comb2ro_0[3:3]);
  OR2 I297 (comb2rro_1[1:1], comb2rr1ltint_0, comb2ro_1[3:3]);
  OR2 I298 (comb2rro_2[1:1], comb2rr1gtint_0, comb2ro_2[3:3]);
  C2 I299 (comb2rro_0[2:2], comb2ro_0[4:4], comb2ro_0[5:5]);
  C2 I300 (comb2rr2ltint_0, comb2ro_1[4:4], comb2ro_0[5:5]);
  C2 I301 (comb2rr2gtint_0, comb2ro_2[4:4], comb2ro_0[5:5]);
  OR2 I302 (comb2rro_1[2:2], comb2rr2ltint_0, comb2ro_1[5:5]);
  OR2 I303 (comb2rro_2[2:2], comb2rr2gtint_0, comb2ro_2[5:5]);
  C2 I304 (comb2rro_0[3:3], comb2ro_0[6:6], comb2ro_0[7:7]);
  C2 I305 (comb2rr3ltint_0, comb2ro_1[6:6], comb2ro_0[7:7]);
  C2 I306 (comb2rr3gtint_0, comb2ro_2[6:6], comb2ro_0[7:7]);
  OR2 I307 (comb2rro_1[3:3], comb2rr3ltint_0, comb2ro_1[7:7]);
  OR2 I308 (comb2rro_2[3:3], comb2rr3gtint_0, comb2ro_2[7:7]);
  C2 I309 (comb2ro_0[0:0], comb2o_0[0:0], comb2o_0[1:1]);
  C2 I310 (comb2r0ltint_0, comb2o_1[0:0], comb2o_0[1:1]);
  C2 I311 (comb2r0gtint_0, comb2o_2[0:0], comb2o_0[1:1]);
  OR2 I312 (comb2ro_1[0:0], comb2r0ltint_0, comb2o_1[1:1]);
  OR2 I313 (comb2ro_2[0:0], comb2r0gtint_0, comb2o_2[1:1]);
  C2 I314 (comb2ro_0[1:1], comb2o_0[2:2], comb2o_0[3:3]);
  C2 I315 (comb2r1ltint_0, comb2o_1[2:2], comb2o_0[3:3]);
  C2 I316 (comb2r1gtint_0, comb2o_2[2:2], comb2o_0[3:3]);
  OR2 I317 (comb2ro_1[1:1], comb2r1ltint_0, comb2o_1[3:3]);
  OR2 I318 (comb2ro_2[1:1], comb2r1gtint_0, comb2o_2[3:3]);
  C2 I319 (comb2ro_0[2:2], comb2o_0[4:4], comb2o_0[5:5]);
  C2 I320 (comb2r2ltint_0, comb2o_1[4:4], comb2o_0[5:5]);
  C2 I321 (comb2r2gtint_0, comb2o_2[4:4], comb2o_0[5:5]);
  OR2 I322 (comb2ro_1[2:2], comb2r2ltint_0, comb2o_1[5:5]);
  OR2 I323 (comb2ro_2[2:2], comb2r2gtint_0, comb2o_2[5:5]);
  C2 I324 (comb2ro_0[3:3], comb2o_0[6:6], comb2o_0[7:7]);
  C2 I325 (comb2r3ltint_0, comb2o_1[6:6], comb2o_0[7:7]);
  C2 I326 (comb2r3gtint_0, comb2o_2[6:6], comb2o_0[7:7]);
  OR2 I327 (comb2ro_1[3:3], comb2r3ltint_0, comb2o_1[7:7]);
  OR2 I328 (comb2ro_2[3:3], comb2r3gtint_0, comb2o_2[7:7]);
  C2 I329 (comb2ro_0[4:4], comb2o_0[8:8], comb2o_0[9:9]);
  C2 I330 (comb2r4ltint_0, comb2o_1[8:8], comb2o_0[9:9]);
  C2 I331 (comb2r4gtint_0, comb2o_2[8:8], comb2o_0[9:9]);
  OR2 I332 (comb2ro_1[4:4], comb2r4ltint_0, comb2o_1[9:9]);
  OR2 I333 (comb2ro_2[4:4], comb2r4gtint_0, comb2o_2[9:9]);
  C2 I334 (comb2ro_0[5:5], comb2o_0[10:10], comb2o_0[11:11]);
  C2 I335 (comb2r5ltint_0, comb2o_1[10:10], comb2o_0[11:11]);
  C2 I336 (comb2r5gtint_0, comb2o_2[10:10], comb2o_0[11:11]);
  OR2 I337 (comb2ro_1[5:5], comb2r5ltint_0, comb2o_1[11:11]);
  OR2 I338 (comb2ro_2[5:5], comb2r5gtint_0, comb2o_2[11:11]);
  C2 I339 (comb2ro_0[6:6], comb2o_0[12:12], comb2o_0[13:13]);
  C2 I340 (comb2r6ltint_0, comb2o_1[12:12], comb2o_0[13:13]);
  C2 I341 (comb2r6gtint_0, comb2o_2[12:12], comb2o_0[13:13]);
  OR2 I342 (comb2ro_1[6:6], comb2r6ltint_0, comb2o_1[13:13]);
  OR2 I343 (comb2ro_2[6:6], comb2r6gtint_0, comb2o_2[13:13]);
  C2 I344 (comb2ro_0[7:7], comb2o_0[14:14], comb2o_0[15:15]);
  C2 I345 (comb2r7ltint_0, comb2o_1[14:14], comb2o_0[15:15]);
  C2 I346 (comb2r7gtint_0, comb2o_2[14:14], comb2o_0[15:15]);
  OR2 I347 (comb2ro_1[7:7], comb2r7ltint_0, comb2o_1[15:15]);
  OR2 I348 (comb2ro_2[7:7], comb2r7gtint_0, comb2o_2[15:15]);
  C2 I349 (comb2o_0[0:0], eq2_0[0:0], eq2_0[1:1]);
  C2 I350 (comb20ltint_0, lt2_0[0:0], eq2_0[1:1]);
  C2 I351 (comb20gtint_0, gt2_0[0:0], eq2_0[1:1]);
  OR2 I352 (comb2o_1[0:0], comb20ltint_0, lt2_0[1:1]);
  OR2 I353 (comb2o_2[0:0], comb20gtint_0, gt2_0[1:1]);
  C2 I354 (comb2o_0[1:1], eq2_0[2:2], eq2_0[3:3]);
  C2 I355 (comb21ltint_0, lt2_0[2:2], eq2_0[3:3]);
  C2 I356 (comb21gtint_0, gt2_0[2:2], eq2_0[3:3]);
  OR2 I357 (comb2o_1[1:1], comb21ltint_0, lt2_0[3:3]);
  OR2 I358 (comb2o_2[1:1], comb21gtint_0, gt2_0[3:3]);
  C2 I359 (comb2o_0[2:2], eq2_0[4:4], eq2_0[5:5]);
  C2 I360 (comb22ltint_0, lt2_0[4:4], eq2_0[5:5]);
  C2 I361 (comb22gtint_0, gt2_0[4:4], eq2_0[5:5]);
  OR2 I362 (comb2o_1[2:2], comb22ltint_0, lt2_0[5:5]);
  OR2 I363 (comb2o_2[2:2], comb22gtint_0, gt2_0[5:5]);
  C2 I364 (comb2o_0[3:3], eq2_0[6:6], eq2_0[7:7]);
  C2 I365 (comb23ltint_0, lt2_0[6:6], eq2_0[7:7]);
  C2 I366 (comb23gtint_0, gt2_0[6:6], eq2_0[7:7]);
  OR2 I367 (comb2o_1[3:3], comb23ltint_0, lt2_0[7:7]);
  OR2 I368 (comb2o_2[3:3], comb23gtint_0, gt2_0[7:7]);
  C2 I369 (comb2o_0[4:4], eq2_0[8:8], eq2_0[9:9]);
  C2 I370 (comb24ltint_0, lt2_0[8:8], eq2_0[9:9]);
  C2 I371 (comb24gtint_0, gt2_0[8:8], eq2_0[9:9]);
  OR2 I372 (comb2o_1[4:4], comb24ltint_0, lt2_0[9:9]);
  OR2 I373 (comb2o_2[4:4], comb24gtint_0, gt2_0[9:9]);
  C2 I374 (comb2o_0[5:5], eq2_0[10:10], eq2_0[11:11]);
  C2 I375 (comb25ltint_0, lt2_0[10:10], eq2_0[11:11]);
  C2 I376 (comb25gtint_0, gt2_0[10:10], eq2_0[11:11]);
  OR2 I377 (comb2o_1[5:5], comb25ltint_0, lt2_0[11:11]);
  OR2 I378 (comb2o_2[5:5], comb25gtint_0, gt2_0[11:11]);
  C2 I379 (comb2o_0[6:6], eq2_0[12:12], eq2_0[13:13]);
  C2 I380 (comb26ltint_0, lt2_0[12:12], eq2_0[13:13]);
  C2 I381 (comb26gtint_0, gt2_0[12:12], eq2_0[13:13]);
  OR2 I382 (comb2o_1[6:6], comb26ltint_0, lt2_0[13:13]);
  OR2 I383 (comb2o_2[6:6], comb26gtint_0, gt2_0[13:13]);
  C2 I384 (comb2o_0[7:7], eq2_0[14:14], eq2_0[15:15]);
  C2 I385 (comb27ltint_0, lt2_0[14:14], eq2_0[15:15]);
  C2 I386 (comb27gtint_0, gt2_0[14:14], eq2_0[15:15]);
  OR2 I387 (comb2o_1[7:7], comb27ltint_0, lt2_0[15:15]);
  OR2 I388 (comb2o_2[7:7], comb27gtint_0, gt2_0[15:15]);
  C2 I389 (comb2o_0[8:8], eq2_0[16:16], eq2_0[17:17]);
  C2 I390 (comb28ltint_0, lt2_0[16:16], eq2_0[17:17]);
  C2 I391 (comb28gtint_0, gt2_0[16:16], eq2_0[17:17]);
  OR2 I392 (comb2o_1[8:8], comb28ltint_0, lt2_0[17:17]);
  OR2 I393 (comb2o_2[8:8], comb28gtint_0, gt2_0[17:17]);
  C2 I394 (comb2o_0[9:9], eq2_0[18:18], eq2_0[19:19]);
  C2 I395 (comb29ltint_0, lt2_0[18:18], eq2_0[19:19]);
  C2 I396 (comb29gtint_0, gt2_0[18:18], eq2_0[19:19]);
  OR2 I397 (comb2o_1[9:9], comb29ltint_0, lt2_0[19:19]);
  OR2 I398 (comb2o_2[9:9], comb29gtint_0, gt2_0[19:19]);
  C2 I399 (comb2o_0[10:10], eq2_0[20:20], eq2_0[21:21]);
  C2 I400 (comb210ltint_0, lt2_0[20:20], eq2_0[21:21]);
  C2 I401 (comb210gtint_0, gt2_0[20:20], eq2_0[21:21]);
  OR2 I402 (comb2o_1[10:10], comb210ltint_0, lt2_0[21:21]);
  OR2 I403 (comb2o_2[10:10], comb210gtint_0, gt2_0[21:21]);
  C2 I404 (comb2o_0[11:11], eq2_0[22:22], eq2_0[23:23]);
  C2 I405 (comb211ltint_0, lt2_0[22:22], eq2_0[23:23]);
  C2 I406 (comb211gtint_0, gt2_0[22:22], eq2_0[23:23]);
  OR2 I407 (comb2o_1[11:11], comb211ltint_0, lt2_0[23:23]);
  OR2 I408 (comb2o_2[11:11], comb211gtint_0, gt2_0[23:23]);
  C2 I409 (comb2o_0[12:12], eq2_0[24:24], eq2_0[25:25]);
  C2 I410 (comb212ltint_0, lt2_0[24:24], eq2_0[25:25]);
  C2 I411 (comb212gtint_0, gt2_0[24:24], eq2_0[25:25]);
  OR2 I412 (comb2o_1[12:12], comb212ltint_0, lt2_0[25:25]);
  OR2 I413 (comb2o_2[12:12], comb212gtint_0, gt2_0[25:25]);
  C2 I414 (comb2o_0[13:13], eq2_0[26:26], eq2_0[27:27]);
  C2 I415 (comb213ltint_0, lt2_0[26:26], eq2_0[27:27]);
  C2 I416 (comb213gtint_0, gt2_0[26:26], eq2_0[27:27]);
  OR2 I417 (comb2o_1[13:13], comb213ltint_0, lt2_0[27:27]);
  OR2 I418 (comb2o_2[13:13], comb213gtint_0, gt2_0[27:27]);
  C2 I419 (comb2o_0[14:14], eq2_0[28:28], eq2_0[29:29]);
  C2 I420 (comb214ltint_0, lt2_0[28:28], eq2_0[29:29]);
  C2 I421 (comb214gtint_0, gt2_0[28:28], eq2_0[29:29]);
  OR2 I422 (comb2o_1[14:14], comb214ltint_0, lt2_0[29:29]);
  OR2 I423 (comb2o_2[14:14], comb214gtint_0, gt2_0[29:29]);
  C2 I424 (comb2o_0[15:15], eq2_0[30:30], eq2_0[31:31]);
  C2 I425 (comb215ltint_0, lt2_0[30:30], eq2_0[31:31]);
  C2 I426 (comb215gtint_0, gt2_0[30:30], eq2_0[31:31]);
  OR2 I427 (comb2o_1[15:15], comb215ltint_0, lt2_0[31:31]);
  OR2 I428 (comb2o_2[15:15], comb215gtint_0, gt2_0[31:31]);
  OR2 I429 (o_0r0, olt2_0, oeq2_0);
  BUFF I430 (o_0r1, ogt2_0);
  BUFF I431 (i_0a, o_0a);
endmodule

// tko32m33_1api0w32bi31w1b_2nm33b1_3subt1o0w33bt2o0w33b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32),(0,31+:1)]),
//     (2,TeakOConstant 33 1),
//     (3,TeakOp TeakOpSub [(1,0+:33),(2,0+:33)])] [One 32,One 33]
module tko32m33_1api0w32bi31w1b_2nm33b1_3subt1o0w33bt2o0w33b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [31:0] gocomp_0;
  wire [10:0] simp341_0;
  wire [3:0] simp342_0;
  wire [1:0] simp343_0;
  wire [32:0] termf_1;
  wire [32:0] termf_2;
  wire [32:0] termt_1;
  wire [32:0] termt_2;
  wire [32:0] cf3__0;
  wire [32:0] ct3__0;
  wire [3:0] ha3__0;
  wire [7:0] fa3_1min_0;
  wire [1:0] simp1291_0;
  wire [1:0] simp1301_0;
  wire [7:0] fa3_2min_0;
  wire [1:0] simp1421_0;
  wire [1:0] simp1431_0;
  wire [7:0] fa3_3min_0;
  wire [1:0] simp1551_0;
  wire [1:0] simp1561_0;
  wire [7:0] fa3_4min_0;
  wire [1:0] simp1681_0;
  wire [1:0] simp1691_0;
  wire [7:0] fa3_5min_0;
  wire [1:0] simp1811_0;
  wire [1:0] simp1821_0;
  wire [7:0] fa3_6min_0;
  wire [1:0] simp1941_0;
  wire [1:0] simp1951_0;
  wire [7:0] fa3_7min_0;
  wire [1:0] simp2071_0;
  wire [1:0] simp2081_0;
  wire [7:0] fa3_8min_0;
  wire [1:0] simp2201_0;
  wire [1:0] simp2211_0;
  wire [7:0] fa3_9min_0;
  wire [1:0] simp2331_0;
  wire [1:0] simp2341_0;
  wire [7:0] fa3_10min_0;
  wire [1:0] simp2461_0;
  wire [1:0] simp2471_0;
  wire [7:0] fa3_11min_0;
  wire [1:0] simp2591_0;
  wire [1:0] simp2601_0;
  wire [7:0] fa3_12min_0;
  wire [1:0] simp2721_0;
  wire [1:0] simp2731_0;
  wire [7:0] fa3_13min_0;
  wire [1:0] simp2851_0;
  wire [1:0] simp2861_0;
  wire [7:0] fa3_14min_0;
  wire [1:0] simp2981_0;
  wire [1:0] simp2991_0;
  wire [7:0] fa3_15min_0;
  wire [1:0] simp3111_0;
  wire [1:0] simp3121_0;
  wire [7:0] fa3_16min_0;
  wire [1:0] simp3241_0;
  wire [1:0] simp3251_0;
  wire [7:0] fa3_17min_0;
  wire [1:0] simp3371_0;
  wire [1:0] simp3381_0;
  wire [7:0] fa3_18min_0;
  wire [1:0] simp3501_0;
  wire [1:0] simp3511_0;
  wire [7:0] fa3_19min_0;
  wire [1:0] simp3631_0;
  wire [1:0] simp3641_0;
  wire [7:0] fa3_20min_0;
  wire [1:0] simp3761_0;
  wire [1:0] simp3771_0;
  wire [7:0] fa3_21min_0;
  wire [1:0] simp3891_0;
  wire [1:0] simp3901_0;
  wire [7:0] fa3_22min_0;
  wire [1:0] simp4021_0;
  wire [1:0] simp4031_0;
  wire [7:0] fa3_23min_0;
  wire [1:0] simp4151_0;
  wire [1:0] simp4161_0;
  wire [7:0] fa3_24min_0;
  wire [1:0] simp4281_0;
  wire [1:0] simp4291_0;
  wire [7:0] fa3_25min_0;
  wire [1:0] simp4411_0;
  wire [1:0] simp4421_0;
  wire [7:0] fa3_26min_0;
  wire [1:0] simp4541_0;
  wire [1:0] simp4551_0;
  wire [7:0] fa3_27min_0;
  wire [1:0] simp4671_0;
  wire [1:0] simp4681_0;
  wire [7:0] fa3_28min_0;
  wire [1:0] simp4801_0;
  wire [1:0] simp4811_0;
  wire [7:0] fa3_29min_0;
  wire [1:0] simp4931_0;
  wire [1:0] simp4941_0;
  wire [7:0] fa3_30min_0;
  wire [1:0] simp5061_0;
  wire [1:0] simp5071_0;
  wire [7:0] fa3_31min_0;
  wire [1:0] simp5191_0;
  wire [1:0] simp5201_0;
  wire [7:0] fa3_32min_0;
  wire [1:0] simp5321_0;
  wire [1:0] simp5331_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I32 (simp341_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I33 (simp341_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I34 (simp341_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I35 (simp341_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I36 (simp341_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I37 (simp341_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I38 (simp341_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I39 (simp341_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I40 (simp341_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I41 (simp341_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C2 I42 (simp341_0[10:10], gocomp_0[30:30], gocomp_0[31:31]);
  C3 I43 (simp342_0[0:0], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  C3 I44 (simp342_0[1:1], simp341_0[3:3], simp341_0[4:4], simp341_0[5:5]);
  C3 I45 (simp342_0[2:2], simp341_0[6:6], simp341_0[7:7], simp341_0[8:8]);
  C2 I46 (simp342_0[3:3], simp341_0[9:9], simp341_0[10:10]);
  C3 I47 (simp343_0[0:0], simp342_0[0:0], simp342_0[1:1], simp342_0[2:2]);
  BUFF I48 (simp343_0[1:1], simp342_0[3:3]);
  C2 I49 (go_0, simp343_0[0:0], simp343_0[1:1]);
  BUFF I50 (termf_1[0:0], i_0r0[0:0]);
  BUFF I51 (termf_1[1:1], i_0r0[1:1]);
  BUFF I52 (termf_1[2:2], i_0r0[2:2]);
  BUFF I53 (termf_1[3:3], i_0r0[3:3]);
  BUFF I54 (termf_1[4:4], i_0r0[4:4]);
  BUFF I55 (termf_1[5:5], i_0r0[5:5]);
  BUFF I56 (termf_1[6:6], i_0r0[6:6]);
  BUFF I57 (termf_1[7:7], i_0r0[7:7]);
  BUFF I58 (termf_1[8:8], i_0r0[8:8]);
  BUFF I59 (termf_1[9:9], i_0r0[9:9]);
  BUFF I60 (termf_1[10:10], i_0r0[10:10]);
  BUFF I61 (termf_1[11:11], i_0r0[11:11]);
  BUFF I62 (termf_1[12:12], i_0r0[12:12]);
  BUFF I63 (termf_1[13:13], i_0r0[13:13]);
  BUFF I64 (termf_1[14:14], i_0r0[14:14]);
  BUFF I65 (termf_1[15:15], i_0r0[15:15]);
  BUFF I66 (termf_1[16:16], i_0r0[16:16]);
  BUFF I67 (termf_1[17:17], i_0r0[17:17]);
  BUFF I68 (termf_1[18:18], i_0r0[18:18]);
  BUFF I69 (termf_1[19:19], i_0r0[19:19]);
  BUFF I70 (termf_1[20:20], i_0r0[20:20]);
  BUFF I71 (termf_1[21:21], i_0r0[21:21]);
  BUFF I72 (termf_1[22:22], i_0r0[22:22]);
  BUFF I73 (termf_1[23:23], i_0r0[23:23]);
  BUFF I74 (termf_1[24:24], i_0r0[24:24]);
  BUFF I75 (termf_1[25:25], i_0r0[25:25]);
  BUFF I76 (termf_1[26:26], i_0r0[26:26]);
  BUFF I77 (termf_1[27:27], i_0r0[27:27]);
  BUFF I78 (termf_1[28:28], i_0r0[28:28]);
  BUFF I79 (termf_1[29:29], i_0r0[29:29]);
  BUFF I80 (termf_1[30:30], i_0r0[30:30]);
  BUFF I81 (termf_1[31:31], i_0r0[31:31]);
  BUFF I82 (termf_1[32:32], i_0r0[31:31]);
  BUFF I83 (termt_1[0:0], i_0r1[0:0]);
  BUFF I84 (termt_1[1:1], i_0r1[1:1]);
  BUFF I85 (termt_1[2:2], i_0r1[2:2]);
  BUFF I86 (termt_1[3:3], i_0r1[3:3]);
  BUFF I87 (termt_1[4:4], i_0r1[4:4]);
  BUFF I88 (termt_1[5:5], i_0r1[5:5]);
  BUFF I89 (termt_1[6:6], i_0r1[6:6]);
  BUFF I90 (termt_1[7:7], i_0r1[7:7]);
  BUFF I91 (termt_1[8:8], i_0r1[8:8]);
  BUFF I92 (termt_1[9:9], i_0r1[9:9]);
  BUFF I93 (termt_1[10:10], i_0r1[10:10]);
  BUFF I94 (termt_1[11:11], i_0r1[11:11]);
  BUFF I95 (termt_1[12:12], i_0r1[12:12]);
  BUFF I96 (termt_1[13:13], i_0r1[13:13]);
  BUFF I97 (termt_1[14:14], i_0r1[14:14]);
  BUFF I98 (termt_1[15:15], i_0r1[15:15]);
  BUFF I99 (termt_1[16:16], i_0r1[16:16]);
  BUFF I100 (termt_1[17:17], i_0r1[17:17]);
  BUFF I101 (termt_1[18:18], i_0r1[18:18]);
  BUFF I102 (termt_1[19:19], i_0r1[19:19]);
  BUFF I103 (termt_1[20:20], i_0r1[20:20]);
  BUFF I104 (termt_1[21:21], i_0r1[21:21]);
  BUFF I105 (termt_1[22:22], i_0r1[22:22]);
  BUFF I106 (termt_1[23:23], i_0r1[23:23]);
  BUFF I107 (termt_1[24:24], i_0r1[24:24]);
  BUFF I108 (termt_1[25:25], i_0r1[25:25]);
  BUFF I109 (termt_1[26:26], i_0r1[26:26]);
  BUFF I110 (termt_1[27:27], i_0r1[27:27]);
  BUFF I111 (termt_1[28:28], i_0r1[28:28]);
  BUFF I112 (termt_1[29:29], i_0r1[29:29]);
  BUFF I113 (termt_1[30:30], i_0r1[30:30]);
  BUFF I114 (termt_1[31:31], i_0r1[31:31]);
  BUFF I115 (termt_1[32:32], i_0r1[31:31]);
  BUFF I116 (termt_2[0:0], go_0);
  GND I117 (termf_2[0:0]);
  BUFF I118 (termf_2[1:1], go_0);
  BUFF I119 (termf_2[2:2], go_0);
  BUFF I120 (termf_2[3:3], go_0);
  BUFF I121 (termf_2[4:4], go_0);
  BUFF I122 (termf_2[5:5], go_0);
  BUFF I123 (termf_2[6:6], go_0);
  BUFF I124 (termf_2[7:7], go_0);
  BUFF I125 (termf_2[8:8], go_0);
  BUFF I126 (termf_2[9:9], go_0);
  BUFF I127 (termf_2[10:10], go_0);
  BUFF I128 (termf_2[11:11], go_0);
  BUFF I129 (termf_2[12:12], go_0);
  BUFF I130 (termf_2[13:13], go_0);
  BUFF I131 (termf_2[14:14], go_0);
  BUFF I132 (termf_2[15:15], go_0);
  BUFF I133 (termf_2[16:16], go_0);
  BUFF I134 (termf_2[17:17], go_0);
  BUFF I135 (termf_2[18:18], go_0);
  BUFF I136 (termf_2[19:19], go_0);
  BUFF I137 (termf_2[20:20], go_0);
  BUFF I138 (termf_2[21:21], go_0);
  BUFF I139 (termf_2[22:22], go_0);
  BUFF I140 (termf_2[23:23], go_0);
  BUFF I141 (termf_2[24:24], go_0);
  BUFF I142 (termf_2[25:25], go_0);
  BUFF I143 (termf_2[26:26], go_0);
  BUFF I144 (termf_2[27:27], go_0);
  BUFF I145 (termf_2[28:28], go_0);
  BUFF I146 (termf_2[29:29], go_0);
  BUFF I147 (termf_2[30:30], go_0);
  BUFF I148 (termf_2[31:31], go_0);
  BUFF I149 (termf_2[32:32], go_0);
  GND I150 (termt_2[1:1]);
  GND I151 (termt_2[2:2]);
  GND I152 (termt_2[3:3]);
  GND I153 (termt_2[4:4]);
  GND I154 (termt_2[5:5]);
  GND I155 (termt_2[6:6]);
  GND I156 (termt_2[7:7]);
  GND I157 (termt_2[8:8]);
  GND I158 (termt_2[9:9]);
  GND I159 (termt_2[10:10]);
  GND I160 (termt_2[11:11]);
  GND I161 (termt_2[12:12]);
  GND I162 (termt_2[13:13]);
  GND I163 (termt_2[14:14]);
  GND I164 (termt_2[15:15]);
  GND I165 (termt_2[16:16]);
  GND I166 (termt_2[17:17]);
  GND I167 (termt_2[18:18]);
  GND I168 (termt_2[19:19]);
  GND I169 (termt_2[20:20]);
  GND I170 (termt_2[21:21]);
  GND I171 (termt_2[22:22]);
  GND I172 (termt_2[23:23]);
  GND I173 (termt_2[24:24]);
  GND I174 (termt_2[25:25]);
  GND I175 (termt_2[26:26]);
  GND I176 (termt_2[27:27]);
  GND I177 (termt_2[28:28]);
  GND I178 (termt_2[29:29]);
  GND I179 (termt_2[30:30]);
  GND I180 (termt_2[31:31]);
  GND I181 (termt_2[32:32]);
  C2 I182 (ha3__0[0:0], termt_2[0:0], termf_1[0:0]);
  C2 I183 (ha3__0[1:1], termt_2[0:0], termt_1[0:0]);
  C2 I184 (ha3__0[2:2], termf_2[0:0], termf_1[0:0]);
  C2 I185 (ha3__0[3:3], termf_2[0:0], termt_1[0:0]);
  BUFF I186 (cf3__0[0:0], ha3__0[0:0]);
  OR3 I187 (ct3__0[0:0], ha3__0[1:1], ha3__0[2:2], ha3__0[3:3]);
  OR2 I188 (o_0r0[0:0], ha3__0[1:1], ha3__0[2:2]);
  OR2 I189 (o_0r1[0:0], ha3__0[0:0], ha3__0[3:3]);
  C3 I190 (fa3_1min_0[0:0], cf3__0[0:0], termt_2[1:1], termf_1[1:1]);
  C3 I191 (fa3_1min_0[1:1], cf3__0[0:0], termt_2[1:1], termt_1[1:1]);
  C3 I192 (fa3_1min_0[2:2], cf3__0[0:0], termf_2[1:1], termf_1[1:1]);
  C3 I193 (fa3_1min_0[3:3], cf3__0[0:0], termf_2[1:1], termt_1[1:1]);
  C3 I194 (fa3_1min_0[4:4], ct3__0[0:0], termt_2[1:1], termf_1[1:1]);
  C3 I195 (fa3_1min_0[5:5], ct3__0[0:0], termt_2[1:1], termt_1[1:1]);
  C3 I196 (fa3_1min_0[6:6], ct3__0[0:0], termf_2[1:1], termf_1[1:1]);
  C3 I197 (fa3_1min_0[7:7], ct3__0[0:0], termf_2[1:1], termt_1[1:1]);
  NOR3 I198 (simp1291_0[0:0], fa3_1min_0[0:0], fa3_1min_0[3:3], fa3_1min_0[5:5]);
  INV I199 (simp1291_0[1:1], fa3_1min_0[6:6]);
  NAND2 I200 (o_0r0[1:1], simp1291_0[0:0], simp1291_0[1:1]);
  NOR3 I201 (simp1301_0[0:0], fa3_1min_0[1:1], fa3_1min_0[2:2], fa3_1min_0[4:4]);
  INV I202 (simp1301_0[1:1], fa3_1min_0[7:7]);
  NAND2 I203 (o_0r1[1:1], simp1301_0[0:0], simp1301_0[1:1]);
  AO222 I204 (ct3__0[1:1], termt_1[1:1], termf_2[1:1], termt_1[1:1], ct3__0[0:0], termf_2[1:1], ct3__0[0:0]);
  AO222 I205 (cf3__0[1:1], termf_1[1:1], termt_2[1:1], termf_1[1:1], cf3__0[0:0], termt_2[1:1], cf3__0[0:0]);
  C3 I206 (fa3_2min_0[0:0], cf3__0[1:1], termt_2[2:2], termf_1[2:2]);
  C3 I207 (fa3_2min_0[1:1], cf3__0[1:1], termt_2[2:2], termt_1[2:2]);
  C3 I208 (fa3_2min_0[2:2], cf3__0[1:1], termf_2[2:2], termf_1[2:2]);
  C3 I209 (fa3_2min_0[3:3], cf3__0[1:1], termf_2[2:2], termt_1[2:2]);
  C3 I210 (fa3_2min_0[4:4], ct3__0[1:1], termt_2[2:2], termf_1[2:2]);
  C3 I211 (fa3_2min_0[5:5], ct3__0[1:1], termt_2[2:2], termt_1[2:2]);
  C3 I212 (fa3_2min_0[6:6], ct3__0[1:1], termf_2[2:2], termf_1[2:2]);
  C3 I213 (fa3_2min_0[7:7], ct3__0[1:1], termf_2[2:2], termt_1[2:2]);
  NOR3 I214 (simp1421_0[0:0], fa3_2min_0[0:0], fa3_2min_0[3:3], fa3_2min_0[5:5]);
  INV I215 (simp1421_0[1:1], fa3_2min_0[6:6]);
  NAND2 I216 (o_0r0[2:2], simp1421_0[0:0], simp1421_0[1:1]);
  NOR3 I217 (simp1431_0[0:0], fa3_2min_0[1:1], fa3_2min_0[2:2], fa3_2min_0[4:4]);
  INV I218 (simp1431_0[1:1], fa3_2min_0[7:7]);
  NAND2 I219 (o_0r1[2:2], simp1431_0[0:0], simp1431_0[1:1]);
  AO222 I220 (ct3__0[2:2], termt_1[2:2], termf_2[2:2], termt_1[2:2], ct3__0[1:1], termf_2[2:2], ct3__0[1:1]);
  AO222 I221 (cf3__0[2:2], termf_1[2:2], termt_2[2:2], termf_1[2:2], cf3__0[1:1], termt_2[2:2], cf3__0[1:1]);
  C3 I222 (fa3_3min_0[0:0], cf3__0[2:2], termt_2[3:3], termf_1[3:3]);
  C3 I223 (fa3_3min_0[1:1], cf3__0[2:2], termt_2[3:3], termt_1[3:3]);
  C3 I224 (fa3_3min_0[2:2], cf3__0[2:2], termf_2[3:3], termf_1[3:3]);
  C3 I225 (fa3_3min_0[3:3], cf3__0[2:2], termf_2[3:3], termt_1[3:3]);
  C3 I226 (fa3_3min_0[4:4], ct3__0[2:2], termt_2[3:3], termf_1[3:3]);
  C3 I227 (fa3_3min_0[5:5], ct3__0[2:2], termt_2[3:3], termt_1[3:3]);
  C3 I228 (fa3_3min_0[6:6], ct3__0[2:2], termf_2[3:3], termf_1[3:3]);
  C3 I229 (fa3_3min_0[7:7], ct3__0[2:2], termf_2[3:3], termt_1[3:3]);
  NOR3 I230 (simp1551_0[0:0], fa3_3min_0[0:0], fa3_3min_0[3:3], fa3_3min_0[5:5]);
  INV I231 (simp1551_0[1:1], fa3_3min_0[6:6]);
  NAND2 I232 (o_0r0[3:3], simp1551_0[0:0], simp1551_0[1:1]);
  NOR3 I233 (simp1561_0[0:0], fa3_3min_0[1:1], fa3_3min_0[2:2], fa3_3min_0[4:4]);
  INV I234 (simp1561_0[1:1], fa3_3min_0[7:7]);
  NAND2 I235 (o_0r1[3:3], simp1561_0[0:0], simp1561_0[1:1]);
  AO222 I236 (ct3__0[3:3], termt_1[3:3], termf_2[3:3], termt_1[3:3], ct3__0[2:2], termf_2[3:3], ct3__0[2:2]);
  AO222 I237 (cf3__0[3:3], termf_1[3:3], termt_2[3:3], termf_1[3:3], cf3__0[2:2], termt_2[3:3], cf3__0[2:2]);
  C3 I238 (fa3_4min_0[0:0], cf3__0[3:3], termt_2[4:4], termf_1[4:4]);
  C3 I239 (fa3_4min_0[1:1], cf3__0[3:3], termt_2[4:4], termt_1[4:4]);
  C3 I240 (fa3_4min_0[2:2], cf3__0[3:3], termf_2[4:4], termf_1[4:4]);
  C3 I241 (fa3_4min_0[3:3], cf3__0[3:3], termf_2[4:4], termt_1[4:4]);
  C3 I242 (fa3_4min_0[4:4], ct3__0[3:3], termt_2[4:4], termf_1[4:4]);
  C3 I243 (fa3_4min_0[5:5], ct3__0[3:3], termt_2[4:4], termt_1[4:4]);
  C3 I244 (fa3_4min_0[6:6], ct3__0[3:3], termf_2[4:4], termf_1[4:4]);
  C3 I245 (fa3_4min_0[7:7], ct3__0[3:3], termf_2[4:4], termt_1[4:4]);
  NOR3 I246 (simp1681_0[0:0], fa3_4min_0[0:0], fa3_4min_0[3:3], fa3_4min_0[5:5]);
  INV I247 (simp1681_0[1:1], fa3_4min_0[6:6]);
  NAND2 I248 (o_0r0[4:4], simp1681_0[0:0], simp1681_0[1:1]);
  NOR3 I249 (simp1691_0[0:0], fa3_4min_0[1:1], fa3_4min_0[2:2], fa3_4min_0[4:4]);
  INV I250 (simp1691_0[1:1], fa3_4min_0[7:7]);
  NAND2 I251 (o_0r1[4:4], simp1691_0[0:0], simp1691_0[1:1]);
  AO222 I252 (ct3__0[4:4], termt_1[4:4], termf_2[4:4], termt_1[4:4], ct3__0[3:3], termf_2[4:4], ct3__0[3:3]);
  AO222 I253 (cf3__0[4:4], termf_1[4:4], termt_2[4:4], termf_1[4:4], cf3__0[3:3], termt_2[4:4], cf3__0[3:3]);
  C3 I254 (fa3_5min_0[0:0], cf3__0[4:4], termt_2[5:5], termf_1[5:5]);
  C3 I255 (fa3_5min_0[1:1], cf3__0[4:4], termt_2[5:5], termt_1[5:5]);
  C3 I256 (fa3_5min_0[2:2], cf3__0[4:4], termf_2[5:5], termf_1[5:5]);
  C3 I257 (fa3_5min_0[3:3], cf3__0[4:4], termf_2[5:5], termt_1[5:5]);
  C3 I258 (fa3_5min_0[4:4], ct3__0[4:4], termt_2[5:5], termf_1[5:5]);
  C3 I259 (fa3_5min_0[5:5], ct3__0[4:4], termt_2[5:5], termt_1[5:5]);
  C3 I260 (fa3_5min_0[6:6], ct3__0[4:4], termf_2[5:5], termf_1[5:5]);
  C3 I261 (fa3_5min_0[7:7], ct3__0[4:4], termf_2[5:5], termt_1[5:5]);
  NOR3 I262 (simp1811_0[0:0], fa3_5min_0[0:0], fa3_5min_0[3:3], fa3_5min_0[5:5]);
  INV I263 (simp1811_0[1:1], fa3_5min_0[6:6]);
  NAND2 I264 (o_0r0[5:5], simp1811_0[0:0], simp1811_0[1:1]);
  NOR3 I265 (simp1821_0[0:0], fa3_5min_0[1:1], fa3_5min_0[2:2], fa3_5min_0[4:4]);
  INV I266 (simp1821_0[1:1], fa3_5min_0[7:7]);
  NAND2 I267 (o_0r1[5:5], simp1821_0[0:0], simp1821_0[1:1]);
  AO222 I268 (ct3__0[5:5], termt_1[5:5], termf_2[5:5], termt_1[5:5], ct3__0[4:4], termf_2[5:5], ct3__0[4:4]);
  AO222 I269 (cf3__0[5:5], termf_1[5:5], termt_2[5:5], termf_1[5:5], cf3__0[4:4], termt_2[5:5], cf3__0[4:4]);
  C3 I270 (fa3_6min_0[0:0], cf3__0[5:5], termt_2[6:6], termf_1[6:6]);
  C3 I271 (fa3_6min_0[1:1], cf3__0[5:5], termt_2[6:6], termt_1[6:6]);
  C3 I272 (fa3_6min_0[2:2], cf3__0[5:5], termf_2[6:6], termf_1[6:6]);
  C3 I273 (fa3_6min_0[3:3], cf3__0[5:5], termf_2[6:6], termt_1[6:6]);
  C3 I274 (fa3_6min_0[4:4], ct3__0[5:5], termt_2[6:6], termf_1[6:6]);
  C3 I275 (fa3_6min_0[5:5], ct3__0[5:5], termt_2[6:6], termt_1[6:6]);
  C3 I276 (fa3_6min_0[6:6], ct3__0[5:5], termf_2[6:6], termf_1[6:6]);
  C3 I277 (fa3_6min_0[7:7], ct3__0[5:5], termf_2[6:6], termt_1[6:6]);
  NOR3 I278 (simp1941_0[0:0], fa3_6min_0[0:0], fa3_6min_0[3:3], fa3_6min_0[5:5]);
  INV I279 (simp1941_0[1:1], fa3_6min_0[6:6]);
  NAND2 I280 (o_0r0[6:6], simp1941_0[0:0], simp1941_0[1:1]);
  NOR3 I281 (simp1951_0[0:0], fa3_6min_0[1:1], fa3_6min_0[2:2], fa3_6min_0[4:4]);
  INV I282 (simp1951_0[1:1], fa3_6min_0[7:7]);
  NAND2 I283 (o_0r1[6:6], simp1951_0[0:0], simp1951_0[1:1]);
  AO222 I284 (ct3__0[6:6], termt_1[6:6], termf_2[6:6], termt_1[6:6], ct3__0[5:5], termf_2[6:6], ct3__0[5:5]);
  AO222 I285 (cf3__0[6:6], termf_1[6:6], termt_2[6:6], termf_1[6:6], cf3__0[5:5], termt_2[6:6], cf3__0[5:5]);
  C3 I286 (fa3_7min_0[0:0], cf3__0[6:6], termt_2[7:7], termf_1[7:7]);
  C3 I287 (fa3_7min_0[1:1], cf3__0[6:6], termt_2[7:7], termt_1[7:7]);
  C3 I288 (fa3_7min_0[2:2], cf3__0[6:6], termf_2[7:7], termf_1[7:7]);
  C3 I289 (fa3_7min_0[3:3], cf3__0[6:6], termf_2[7:7], termt_1[7:7]);
  C3 I290 (fa3_7min_0[4:4], ct3__0[6:6], termt_2[7:7], termf_1[7:7]);
  C3 I291 (fa3_7min_0[5:5], ct3__0[6:6], termt_2[7:7], termt_1[7:7]);
  C3 I292 (fa3_7min_0[6:6], ct3__0[6:6], termf_2[7:7], termf_1[7:7]);
  C3 I293 (fa3_7min_0[7:7], ct3__0[6:6], termf_2[7:7], termt_1[7:7]);
  NOR3 I294 (simp2071_0[0:0], fa3_7min_0[0:0], fa3_7min_0[3:3], fa3_7min_0[5:5]);
  INV I295 (simp2071_0[1:1], fa3_7min_0[6:6]);
  NAND2 I296 (o_0r0[7:7], simp2071_0[0:0], simp2071_0[1:1]);
  NOR3 I297 (simp2081_0[0:0], fa3_7min_0[1:1], fa3_7min_0[2:2], fa3_7min_0[4:4]);
  INV I298 (simp2081_0[1:1], fa3_7min_0[7:7]);
  NAND2 I299 (o_0r1[7:7], simp2081_0[0:0], simp2081_0[1:1]);
  AO222 I300 (ct3__0[7:7], termt_1[7:7], termf_2[7:7], termt_1[7:7], ct3__0[6:6], termf_2[7:7], ct3__0[6:6]);
  AO222 I301 (cf3__0[7:7], termf_1[7:7], termt_2[7:7], termf_1[7:7], cf3__0[6:6], termt_2[7:7], cf3__0[6:6]);
  C3 I302 (fa3_8min_0[0:0], cf3__0[7:7], termt_2[8:8], termf_1[8:8]);
  C3 I303 (fa3_8min_0[1:1], cf3__0[7:7], termt_2[8:8], termt_1[8:8]);
  C3 I304 (fa3_8min_0[2:2], cf3__0[7:7], termf_2[8:8], termf_1[8:8]);
  C3 I305 (fa3_8min_0[3:3], cf3__0[7:7], termf_2[8:8], termt_1[8:8]);
  C3 I306 (fa3_8min_0[4:4], ct3__0[7:7], termt_2[8:8], termf_1[8:8]);
  C3 I307 (fa3_8min_0[5:5], ct3__0[7:7], termt_2[8:8], termt_1[8:8]);
  C3 I308 (fa3_8min_0[6:6], ct3__0[7:7], termf_2[8:8], termf_1[8:8]);
  C3 I309 (fa3_8min_0[7:7], ct3__0[7:7], termf_2[8:8], termt_1[8:8]);
  NOR3 I310 (simp2201_0[0:0], fa3_8min_0[0:0], fa3_8min_0[3:3], fa3_8min_0[5:5]);
  INV I311 (simp2201_0[1:1], fa3_8min_0[6:6]);
  NAND2 I312 (o_0r0[8:8], simp2201_0[0:0], simp2201_0[1:1]);
  NOR3 I313 (simp2211_0[0:0], fa3_8min_0[1:1], fa3_8min_0[2:2], fa3_8min_0[4:4]);
  INV I314 (simp2211_0[1:1], fa3_8min_0[7:7]);
  NAND2 I315 (o_0r1[8:8], simp2211_0[0:0], simp2211_0[1:1]);
  AO222 I316 (ct3__0[8:8], termt_1[8:8], termf_2[8:8], termt_1[8:8], ct3__0[7:7], termf_2[8:8], ct3__0[7:7]);
  AO222 I317 (cf3__0[8:8], termf_1[8:8], termt_2[8:8], termf_1[8:8], cf3__0[7:7], termt_2[8:8], cf3__0[7:7]);
  C3 I318 (fa3_9min_0[0:0], cf3__0[8:8], termt_2[9:9], termf_1[9:9]);
  C3 I319 (fa3_9min_0[1:1], cf3__0[8:8], termt_2[9:9], termt_1[9:9]);
  C3 I320 (fa3_9min_0[2:2], cf3__0[8:8], termf_2[9:9], termf_1[9:9]);
  C3 I321 (fa3_9min_0[3:3], cf3__0[8:8], termf_2[9:9], termt_1[9:9]);
  C3 I322 (fa3_9min_0[4:4], ct3__0[8:8], termt_2[9:9], termf_1[9:9]);
  C3 I323 (fa3_9min_0[5:5], ct3__0[8:8], termt_2[9:9], termt_1[9:9]);
  C3 I324 (fa3_9min_0[6:6], ct3__0[8:8], termf_2[9:9], termf_1[9:9]);
  C3 I325 (fa3_9min_0[7:7], ct3__0[8:8], termf_2[9:9], termt_1[9:9]);
  NOR3 I326 (simp2331_0[0:0], fa3_9min_0[0:0], fa3_9min_0[3:3], fa3_9min_0[5:5]);
  INV I327 (simp2331_0[1:1], fa3_9min_0[6:6]);
  NAND2 I328 (o_0r0[9:9], simp2331_0[0:0], simp2331_0[1:1]);
  NOR3 I329 (simp2341_0[0:0], fa3_9min_0[1:1], fa3_9min_0[2:2], fa3_9min_0[4:4]);
  INV I330 (simp2341_0[1:1], fa3_9min_0[7:7]);
  NAND2 I331 (o_0r1[9:9], simp2341_0[0:0], simp2341_0[1:1]);
  AO222 I332 (ct3__0[9:9], termt_1[9:9], termf_2[9:9], termt_1[9:9], ct3__0[8:8], termf_2[9:9], ct3__0[8:8]);
  AO222 I333 (cf3__0[9:9], termf_1[9:9], termt_2[9:9], termf_1[9:9], cf3__0[8:8], termt_2[9:9], cf3__0[8:8]);
  C3 I334 (fa3_10min_0[0:0], cf3__0[9:9], termt_2[10:10], termf_1[10:10]);
  C3 I335 (fa3_10min_0[1:1], cf3__0[9:9], termt_2[10:10], termt_1[10:10]);
  C3 I336 (fa3_10min_0[2:2], cf3__0[9:9], termf_2[10:10], termf_1[10:10]);
  C3 I337 (fa3_10min_0[3:3], cf3__0[9:9], termf_2[10:10], termt_1[10:10]);
  C3 I338 (fa3_10min_0[4:4], ct3__0[9:9], termt_2[10:10], termf_1[10:10]);
  C3 I339 (fa3_10min_0[5:5], ct3__0[9:9], termt_2[10:10], termt_1[10:10]);
  C3 I340 (fa3_10min_0[6:6], ct3__0[9:9], termf_2[10:10], termf_1[10:10]);
  C3 I341 (fa3_10min_0[7:7], ct3__0[9:9], termf_2[10:10], termt_1[10:10]);
  NOR3 I342 (simp2461_0[0:0], fa3_10min_0[0:0], fa3_10min_0[3:3], fa3_10min_0[5:5]);
  INV I343 (simp2461_0[1:1], fa3_10min_0[6:6]);
  NAND2 I344 (o_0r0[10:10], simp2461_0[0:0], simp2461_0[1:1]);
  NOR3 I345 (simp2471_0[0:0], fa3_10min_0[1:1], fa3_10min_0[2:2], fa3_10min_0[4:4]);
  INV I346 (simp2471_0[1:1], fa3_10min_0[7:7]);
  NAND2 I347 (o_0r1[10:10], simp2471_0[0:0], simp2471_0[1:1]);
  AO222 I348 (ct3__0[10:10], termt_1[10:10], termf_2[10:10], termt_1[10:10], ct3__0[9:9], termf_2[10:10], ct3__0[9:9]);
  AO222 I349 (cf3__0[10:10], termf_1[10:10], termt_2[10:10], termf_1[10:10], cf3__0[9:9], termt_2[10:10], cf3__0[9:9]);
  C3 I350 (fa3_11min_0[0:0], cf3__0[10:10], termt_2[11:11], termf_1[11:11]);
  C3 I351 (fa3_11min_0[1:1], cf3__0[10:10], termt_2[11:11], termt_1[11:11]);
  C3 I352 (fa3_11min_0[2:2], cf3__0[10:10], termf_2[11:11], termf_1[11:11]);
  C3 I353 (fa3_11min_0[3:3], cf3__0[10:10], termf_2[11:11], termt_1[11:11]);
  C3 I354 (fa3_11min_0[4:4], ct3__0[10:10], termt_2[11:11], termf_1[11:11]);
  C3 I355 (fa3_11min_0[5:5], ct3__0[10:10], termt_2[11:11], termt_1[11:11]);
  C3 I356 (fa3_11min_0[6:6], ct3__0[10:10], termf_2[11:11], termf_1[11:11]);
  C3 I357 (fa3_11min_0[7:7], ct3__0[10:10], termf_2[11:11], termt_1[11:11]);
  NOR3 I358 (simp2591_0[0:0], fa3_11min_0[0:0], fa3_11min_0[3:3], fa3_11min_0[5:5]);
  INV I359 (simp2591_0[1:1], fa3_11min_0[6:6]);
  NAND2 I360 (o_0r0[11:11], simp2591_0[0:0], simp2591_0[1:1]);
  NOR3 I361 (simp2601_0[0:0], fa3_11min_0[1:1], fa3_11min_0[2:2], fa3_11min_0[4:4]);
  INV I362 (simp2601_0[1:1], fa3_11min_0[7:7]);
  NAND2 I363 (o_0r1[11:11], simp2601_0[0:0], simp2601_0[1:1]);
  AO222 I364 (ct3__0[11:11], termt_1[11:11], termf_2[11:11], termt_1[11:11], ct3__0[10:10], termf_2[11:11], ct3__0[10:10]);
  AO222 I365 (cf3__0[11:11], termf_1[11:11], termt_2[11:11], termf_1[11:11], cf3__0[10:10], termt_2[11:11], cf3__0[10:10]);
  C3 I366 (fa3_12min_0[0:0], cf3__0[11:11], termt_2[12:12], termf_1[12:12]);
  C3 I367 (fa3_12min_0[1:1], cf3__0[11:11], termt_2[12:12], termt_1[12:12]);
  C3 I368 (fa3_12min_0[2:2], cf3__0[11:11], termf_2[12:12], termf_1[12:12]);
  C3 I369 (fa3_12min_0[3:3], cf3__0[11:11], termf_2[12:12], termt_1[12:12]);
  C3 I370 (fa3_12min_0[4:4], ct3__0[11:11], termt_2[12:12], termf_1[12:12]);
  C3 I371 (fa3_12min_0[5:5], ct3__0[11:11], termt_2[12:12], termt_1[12:12]);
  C3 I372 (fa3_12min_0[6:6], ct3__0[11:11], termf_2[12:12], termf_1[12:12]);
  C3 I373 (fa3_12min_0[7:7], ct3__0[11:11], termf_2[12:12], termt_1[12:12]);
  NOR3 I374 (simp2721_0[0:0], fa3_12min_0[0:0], fa3_12min_0[3:3], fa3_12min_0[5:5]);
  INV I375 (simp2721_0[1:1], fa3_12min_0[6:6]);
  NAND2 I376 (o_0r0[12:12], simp2721_0[0:0], simp2721_0[1:1]);
  NOR3 I377 (simp2731_0[0:0], fa3_12min_0[1:1], fa3_12min_0[2:2], fa3_12min_0[4:4]);
  INV I378 (simp2731_0[1:1], fa3_12min_0[7:7]);
  NAND2 I379 (o_0r1[12:12], simp2731_0[0:0], simp2731_0[1:1]);
  AO222 I380 (ct3__0[12:12], termt_1[12:12], termf_2[12:12], termt_1[12:12], ct3__0[11:11], termf_2[12:12], ct3__0[11:11]);
  AO222 I381 (cf3__0[12:12], termf_1[12:12], termt_2[12:12], termf_1[12:12], cf3__0[11:11], termt_2[12:12], cf3__0[11:11]);
  C3 I382 (fa3_13min_0[0:0], cf3__0[12:12], termt_2[13:13], termf_1[13:13]);
  C3 I383 (fa3_13min_0[1:1], cf3__0[12:12], termt_2[13:13], termt_1[13:13]);
  C3 I384 (fa3_13min_0[2:2], cf3__0[12:12], termf_2[13:13], termf_1[13:13]);
  C3 I385 (fa3_13min_0[3:3], cf3__0[12:12], termf_2[13:13], termt_1[13:13]);
  C3 I386 (fa3_13min_0[4:4], ct3__0[12:12], termt_2[13:13], termf_1[13:13]);
  C3 I387 (fa3_13min_0[5:5], ct3__0[12:12], termt_2[13:13], termt_1[13:13]);
  C3 I388 (fa3_13min_0[6:6], ct3__0[12:12], termf_2[13:13], termf_1[13:13]);
  C3 I389 (fa3_13min_0[7:7], ct3__0[12:12], termf_2[13:13], termt_1[13:13]);
  NOR3 I390 (simp2851_0[0:0], fa3_13min_0[0:0], fa3_13min_0[3:3], fa3_13min_0[5:5]);
  INV I391 (simp2851_0[1:1], fa3_13min_0[6:6]);
  NAND2 I392 (o_0r0[13:13], simp2851_0[0:0], simp2851_0[1:1]);
  NOR3 I393 (simp2861_0[0:0], fa3_13min_0[1:1], fa3_13min_0[2:2], fa3_13min_0[4:4]);
  INV I394 (simp2861_0[1:1], fa3_13min_0[7:7]);
  NAND2 I395 (o_0r1[13:13], simp2861_0[0:0], simp2861_0[1:1]);
  AO222 I396 (ct3__0[13:13], termt_1[13:13], termf_2[13:13], termt_1[13:13], ct3__0[12:12], termf_2[13:13], ct3__0[12:12]);
  AO222 I397 (cf3__0[13:13], termf_1[13:13], termt_2[13:13], termf_1[13:13], cf3__0[12:12], termt_2[13:13], cf3__0[12:12]);
  C3 I398 (fa3_14min_0[0:0], cf3__0[13:13], termt_2[14:14], termf_1[14:14]);
  C3 I399 (fa3_14min_0[1:1], cf3__0[13:13], termt_2[14:14], termt_1[14:14]);
  C3 I400 (fa3_14min_0[2:2], cf3__0[13:13], termf_2[14:14], termf_1[14:14]);
  C3 I401 (fa3_14min_0[3:3], cf3__0[13:13], termf_2[14:14], termt_1[14:14]);
  C3 I402 (fa3_14min_0[4:4], ct3__0[13:13], termt_2[14:14], termf_1[14:14]);
  C3 I403 (fa3_14min_0[5:5], ct3__0[13:13], termt_2[14:14], termt_1[14:14]);
  C3 I404 (fa3_14min_0[6:6], ct3__0[13:13], termf_2[14:14], termf_1[14:14]);
  C3 I405 (fa3_14min_0[7:7], ct3__0[13:13], termf_2[14:14], termt_1[14:14]);
  NOR3 I406 (simp2981_0[0:0], fa3_14min_0[0:0], fa3_14min_0[3:3], fa3_14min_0[5:5]);
  INV I407 (simp2981_0[1:1], fa3_14min_0[6:6]);
  NAND2 I408 (o_0r0[14:14], simp2981_0[0:0], simp2981_0[1:1]);
  NOR3 I409 (simp2991_0[0:0], fa3_14min_0[1:1], fa3_14min_0[2:2], fa3_14min_0[4:4]);
  INV I410 (simp2991_0[1:1], fa3_14min_0[7:7]);
  NAND2 I411 (o_0r1[14:14], simp2991_0[0:0], simp2991_0[1:1]);
  AO222 I412 (ct3__0[14:14], termt_1[14:14], termf_2[14:14], termt_1[14:14], ct3__0[13:13], termf_2[14:14], ct3__0[13:13]);
  AO222 I413 (cf3__0[14:14], termf_1[14:14], termt_2[14:14], termf_1[14:14], cf3__0[13:13], termt_2[14:14], cf3__0[13:13]);
  C3 I414 (fa3_15min_0[0:0], cf3__0[14:14], termt_2[15:15], termf_1[15:15]);
  C3 I415 (fa3_15min_0[1:1], cf3__0[14:14], termt_2[15:15], termt_1[15:15]);
  C3 I416 (fa3_15min_0[2:2], cf3__0[14:14], termf_2[15:15], termf_1[15:15]);
  C3 I417 (fa3_15min_0[3:3], cf3__0[14:14], termf_2[15:15], termt_1[15:15]);
  C3 I418 (fa3_15min_0[4:4], ct3__0[14:14], termt_2[15:15], termf_1[15:15]);
  C3 I419 (fa3_15min_0[5:5], ct3__0[14:14], termt_2[15:15], termt_1[15:15]);
  C3 I420 (fa3_15min_0[6:6], ct3__0[14:14], termf_2[15:15], termf_1[15:15]);
  C3 I421 (fa3_15min_0[7:7], ct3__0[14:14], termf_2[15:15], termt_1[15:15]);
  NOR3 I422 (simp3111_0[0:0], fa3_15min_0[0:0], fa3_15min_0[3:3], fa3_15min_0[5:5]);
  INV I423 (simp3111_0[1:1], fa3_15min_0[6:6]);
  NAND2 I424 (o_0r0[15:15], simp3111_0[0:0], simp3111_0[1:1]);
  NOR3 I425 (simp3121_0[0:0], fa3_15min_0[1:1], fa3_15min_0[2:2], fa3_15min_0[4:4]);
  INV I426 (simp3121_0[1:1], fa3_15min_0[7:7]);
  NAND2 I427 (o_0r1[15:15], simp3121_0[0:0], simp3121_0[1:1]);
  AO222 I428 (ct3__0[15:15], termt_1[15:15], termf_2[15:15], termt_1[15:15], ct3__0[14:14], termf_2[15:15], ct3__0[14:14]);
  AO222 I429 (cf3__0[15:15], termf_1[15:15], termt_2[15:15], termf_1[15:15], cf3__0[14:14], termt_2[15:15], cf3__0[14:14]);
  C3 I430 (fa3_16min_0[0:0], cf3__0[15:15], termt_2[16:16], termf_1[16:16]);
  C3 I431 (fa3_16min_0[1:1], cf3__0[15:15], termt_2[16:16], termt_1[16:16]);
  C3 I432 (fa3_16min_0[2:2], cf3__0[15:15], termf_2[16:16], termf_1[16:16]);
  C3 I433 (fa3_16min_0[3:3], cf3__0[15:15], termf_2[16:16], termt_1[16:16]);
  C3 I434 (fa3_16min_0[4:4], ct3__0[15:15], termt_2[16:16], termf_1[16:16]);
  C3 I435 (fa3_16min_0[5:5], ct3__0[15:15], termt_2[16:16], termt_1[16:16]);
  C3 I436 (fa3_16min_0[6:6], ct3__0[15:15], termf_2[16:16], termf_1[16:16]);
  C3 I437 (fa3_16min_0[7:7], ct3__0[15:15], termf_2[16:16], termt_1[16:16]);
  NOR3 I438 (simp3241_0[0:0], fa3_16min_0[0:0], fa3_16min_0[3:3], fa3_16min_0[5:5]);
  INV I439 (simp3241_0[1:1], fa3_16min_0[6:6]);
  NAND2 I440 (o_0r0[16:16], simp3241_0[0:0], simp3241_0[1:1]);
  NOR3 I441 (simp3251_0[0:0], fa3_16min_0[1:1], fa3_16min_0[2:2], fa3_16min_0[4:4]);
  INV I442 (simp3251_0[1:1], fa3_16min_0[7:7]);
  NAND2 I443 (o_0r1[16:16], simp3251_0[0:0], simp3251_0[1:1]);
  AO222 I444 (ct3__0[16:16], termt_1[16:16], termf_2[16:16], termt_1[16:16], ct3__0[15:15], termf_2[16:16], ct3__0[15:15]);
  AO222 I445 (cf3__0[16:16], termf_1[16:16], termt_2[16:16], termf_1[16:16], cf3__0[15:15], termt_2[16:16], cf3__0[15:15]);
  C3 I446 (fa3_17min_0[0:0], cf3__0[16:16], termt_2[17:17], termf_1[17:17]);
  C3 I447 (fa3_17min_0[1:1], cf3__0[16:16], termt_2[17:17], termt_1[17:17]);
  C3 I448 (fa3_17min_0[2:2], cf3__0[16:16], termf_2[17:17], termf_1[17:17]);
  C3 I449 (fa3_17min_0[3:3], cf3__0[16:16], termf_2[17:17], termt_1[17:17]);
  C3 I450 (fa3_17min_0[4:4], ct3__0[16:16], termt_2[17:17], termf_1[17:17]);
  C3 I451 (fa3_17min_0[5:5], ct3__0[16:16], termt_2[17:17], termt_1[17:17]);
  C3 I452 (fa3_17min_0[6:6], ct3__0[16:16], termf_2[17:17], termf_1[17:17]);
  C3 I453 (fa3_17min_0[7:7], ct3__0[16:16], termf_2[17:17], termt_1[17:17]);
  NOR3 I454 (simp3371_0[0:0], fa3_17min_0[0:0], fa3_17min_0[3:3], fa3_17min_0[5:5]);
  INV I455 (simp3371_0[1:1], fa3_17min_0[6:6]);
  NAND2 I456 (o_0r0[17:17], simp3371_0[0:0], simp3371_0[1:1]);
  NOR3 I457 (simp3381_0[0:0], fa3_17min_0[1:1], fa3_17min_0[2:2], fa3_17min_0[4:4]);
  INV I458 (simp3381_0[1:1], fa3_17min_0[7:7]);
  NAND2 I459 (o_0r1[17:17], simp3381_0[0:0], simp3381_0[1:1]);
  AO222 I460 (ct3__0[17:17], termt_1[17:17], termf_2[17:17], termt_1[17:17], ct3__0[16:16], termf_2[17:17], ct3__0[16:16]);
  AO222 I461 (cf3__0[17:17], termf_1[17:17], termt_2[17:17], termf_1[17:17], cf3__0[16:16], termt_2[17:17], cf3__0[16:16]);
  C3 I462 (fa3_18min_0[0:0], cf3__0[17:17], termt_2[18:18], termf_1[18:18]);
  C3 I463 (fa3_18min_0[1:1], cf3__0[17:17], termt_2[18:18], termt_1[18:18]);
  C3 I464 (fa3_18min_0[2:2], cf3__0[17:17], termf_2[18:18], termf_1[18:18]);
  C3 I465 (fa3_18min_0[3:3], cf3__0[17:17], termf_2[18:18], termt_1[18:18]);
  C3 I466 (fa3_18min_0[4:4], ct3__0[17:17], termt_2[18:18], termf_1[18:18]);
  C3 I467 (fa3_18min_0[5:5], ct3__0[17:17], termt_2[18:18], termt_1[18:18]);
  C3 I468 (fa3_18min_0[6:6], ct3__0[17:17], termf_2[18:18], termf_1[18:18]);
  C3 I469 (fa3_18min_0[7:7], ct3__0[17:17], termf_2[18:18], termt_1[18:18]);
  NOR3 I470 (simp3501_0[0:0], fa3_18min_0[0:0], fa3_18min_0[3:3], fa3_18min_0[5:5]);
  INV I471 (simp3501_0[1:1], fa3_18min_0[6:6]);
  NAND2 I472 (o_0r0[18:18], simp3501_0[0:0], simp3501_0[1:1]);
  NOR3 I473 (simp3511_0[0:0], fa3_18min_0[1:1], fa3_18min_0[2:2], fa3_18min_0[4:4]);
  INV I474 (simp3511_0[1:1], fa3_18min_0[7:7]);
  NAND2 I475 (o_0r1[18:18], simp3511_0[0:0], simp3511_0[1:1]);
  AO222 I476 (ct3__0[18:18], termt_1[18:18], termf_2[18:18], termt_1[18:18], ct3__0[17:17], termf_2[18:18], ct3__0[17:17]);
  AO222 I477 (cf3__0[18:18], termf_1[18:18], termt_2[18:18], termf_1[18:18], cf3__0[17:17], termt_2[18:18], cf3__0[17:17]);
  C3 I478 (fa3_19min_0[0:0], cf3__0[18:18], termt_2[19:19], termf_1[19:19]);
  C3 I479 (fa3_19min_0[1:1], cf3__0[18:18], termt_2[19:19], termt_1[19:19]);
  C3 I480 (fa3_19min_0[2:2], cf3__0[18:18], termf_2[19:19], termf_1[19:19]);
  C3 I481 (fa3_19min_0[3:3], cf3__0[18:18], termf_2[19:19], termt_1[19:19]);
  C3 I482 (fa3_19min_0[4:4], ct3__0[18:18], termt_2[19:19], termf_1[19:19]);
  C3 I483 (fa3_19min_0[5:5], ct3__0[18:18], termt_2[19:19], termt_1[19:19]);
  C3 I484 (fa3_19min_0[6:6], ct3__0[18:18], termf_2[19:19], termf_1[19:19]);
  C3 I485 (fa3_19min_0[7:7], ct3__0[18:18], termf_2[19:19], termt_1[19:19]);
  NOR3 I486 (simp3631_0[0:0], fa3_19min_0[0:0], fa3_19min_0[3:3], fa3_19min_0[5:5]);
  INV I487 (simp3631_0[1:1], fa3_19min_0[6:6]);
  NAND2 I488 (o_0r0[19:19], simp3631_0[0:0], simp3631_0[1:1]);
  NOR3 I489 (simp3641_0[0:0], fa3_19min_0[1:1], fa3_19min_0[2:2], fa3_19min_0[4:4]);
  INV I490 (simp3641_0[1:1], fa3_19min_0[7:7]);
  NAND2 I491 (o_0r1[19:19], simp3641_0[0:0], simp3641_0[1:1]);
  AO222 I492 (ct3__0[19:19], termt_1[19:19], termf_2[19:19], termt_1[19:19], ct3__0[18:18], termf_2[19:19], ct3__0[18:18]);
  AO222 I493 (cf3__0[19:19], termf_1[19:19], termt_2[19:19], termf_1[19:19], cf3__0[18:18], termt_2[19:19], cf3__0[18:18]);
  C3 I494 (fa3_20min_0[0:0], cf3__0[19:19], termt_2[20:20], termf_1[20:20]);
  C3 I495 (fa3_20min_0[1:1], cf3__0[19:19], termt_2[20:20], termt_1[20:20]);
  C3 I496 (fa3_20min_0[2:2], cf3__0[19:19], termf_2[20:20], termf_1[20:20]);
  C3 I497 (fa3_20min_0[3:3], cf3__0[19:19], termf_2[20:20], termt_1[20:20]);
  C3 I498 (fa3_20min_0[4:4], ct3__0[19:19], termt_2[20:20], termf_1[20:20]);
  C3 I499 (fa3_20min_0[5:5], ct3__0[19:19], termt_2[20:20], termt_1[20:20]);
  C3 I500 (fa3_20min_0[6:6], ct3__0[19:19], termf_2[20:20], termf_1[20:20]);
  C3 I501 (fa3_20min_0[7:7], ct3__0[19:19], termf_2[20:20], termt_1[20:20]);
  NOR3 I502 (simp3761_0[0:0], fa3_20min_0[0:0], fa3_20min_0[3:3], fa3_20min_0[5:5]);
  INV I503 (simp3761_0[1:1], fa3_20min_0[6:6]);
  NAND2 I504 (o_0r0[20:20], simp3761_0[0:0], simp3761_0[1:1]);
  NOR3 I505 (simp3771_0[0:0], fa3_20min_0[1:1], fa3_20min_0[2:2], fa3_20min_0[4:4]);
  INV I506 (simp3771_0[1:1], fa3_20min_0[7:7]);
  NAND2 I507 (o_0r1[20:20], simp3771_0[0:0], simp3771_0[1:1]);
  AO222 I508 (ct3__0[20:20], termt_1[20:20], termf_2[20:20], termt_1[20:20], ct3__0[19:19], termf_2[20:20], ct3__0[19:19]);
  AO222 I509 (cf3__0[20:20], termf_1[20:20], termt_2[20:20], termf_1[20:20], cf3__0[19:19], termt_2[20:20], cf3__0[19:19]);
  C3 I510 (fa3_21min_0[0:0], cf3__0[20:20], termt_2[21:21], termf_1[21:21]);
  C3 I511 (fa3_21min_0[1:1], cf3__0[20:20], termt_2[21:21], termt_1[21:21]);
  C3 I512 (fa3_21min_0[2:2], cf3__0[20:20], termf_2[21:21], termf_1[21:21]);
  C3 I513 (fa3_21min_0[3:3], cf3__0[20:20], termf_2[21:21], termt_1[21:21]);
  C3 I514 (fa3_21min_0[4:4], ct3__0[20:20], termt_2[21:21], termf_1[21:21]);
  C3 I515 (fa3_21min_0[5:5], ct3__0[20:20], termt_2[21:21], termt_1[21:21]);
  C3 I516 (fa3_21min_0[6:6], ct3__0[20:20], termf_2[21:21], termf_1[21:21]);
  C3 I517 (fa3_21min_0[7:7], ct3__0[20:20], termf_2[21:21], termt_1[21:21]);
  NOR3 I518 (simp3891_0[0:0], fa3_21min_0[0:0], fa3_21min_0[3:3], fa3_21min_0[5:5]);
  INV I519 (simp3891_0[1:1], fa3_21min_0[6:6]);
  NAND2 I520 (o_0r0[21:21], simp3891_0[0:0], simp3891_0[1:1]);
  NOR3 I521 (simp3901_0[0:0], fa3_21min_0[1:1], fa3_21min_0[2:2], fa3_21min_0[4:4]);
  INV I522 (simp3901_0[1:1], fa3_21min_0[7:7]);
  NAND2 I523 (o_0r1[21:21], simp3901_0[0:0], simp3901_0[1:1]);
  AO222 I524 (ct3__0[21:21], termt_1[21:21], termf_2[21:21], termt_1[21:21], ct3__0[20:20], termf_2[21:21], ct3__0[20:20]);
  AO222 I525 (cf3__0[21:21], termf_1[21:21], termt_2[21:21], termf_1[21:21], cf3__0[20:20], termt_2[21:21], cf3__0[20:20]);
  C3 I526 (fa3_22min_0[0:0], cf3__0[21:21], termt_2[22:22], termf_1[22:22]);
  C3 I527 (fa3_22min_0[1:1], cf3__0[21:21], termt_2[22:22], termt_1[22:22]);
  C3 I528 (fa3_22min_0[2:2], cf3__0[21:21], termf_2[22:22], termf_1[22:22]);
  C3 I529 (fa3_22min_0[3:3], cf3__0[21:21], termf_2[22:22], termt_1[22:22]);
  C3 I530 (fa3_22min_0[4:4], ct3__0[21:21], termt_2[22:22], termf_1[22:22]);
  C3 I531 (fa3_22min_0[5:5], ct3__0[21:21], termt_2[22:22], termt_1[22:22]);
  C3 I532 (fa3_22min_0[6:6], ct3__0[21:21], termf_2[22:22], termf_1[22:22]);
  C3 I533 (fa3_22min_0[7:7], ct3__0[21:21], termf_2[22:22], termt_1[22:22]);
  NOR3 I534 (simp4021_0[0:0], fa3_22min_0[0:0], fa3_22min_0[3:3], fa3_22min_0[5:5]);
  INV I535 (simp4021_0[1:1], fa3_22min_0[6:6]);
  NAND2 I536 (o_0r0[22:22], simp4021_0[0:0], simp4021_0[1:1]);
  NOR3 I537 (simp4031_0[0:0], fa3_22min_0[1:1], fa3_22min_0[2:2], fa3_22min_0[4:4]);
  INV I538 (simp4031_0[1:1], fa3_22min_0[7:7]);
  NAND2 I539 (o_0r1[22:22], simp4031_0[0:0], simp4031_0[1:1]);
  AO222 I540 (ct3__0[22:22], termt_1[22:22], termf_2[22:22], termt_1[22:22], ct3__0[21:21], termf_2[22:22], ct3__0[21:21]);
  AO222 I541 (cf3__0[22:22], termf_1[22:22], termt_2[22:22], termf_1[22:22], cf3__0[21:21], termt_2[22:22], cf3__0[21:21]);
  C3 I542 (fa3_23min_0[0:0], cf3__0[22:22], termt_2[23:23], termf_1[23:23]);
  C3 I543 (fa3_23min_0[1:1], cf3__0[22:22], termt_2[23:23], termt_1[23:23]);
  C3 I544 (fa3_23min_0[2:2], cf3__0[22:22], termf_2[23:23], termf_1[23:23]);
  C3 I545 (fa3_23min_0[3:3], cf3__0[22:22], termf_2[23:23], termt_1[23:23]);
  C3 I546 (fa3_23min_0[4:4], ct3__0[22:22], termt_2[23:23], termf_1[23:23]);
  C3 I547 (fa3_23min_0[5:5], ct3__0[22:22], termt_2[23:23], termt_1[23:23]);
  C3 I548 (fa3_23min_0[6:6], ct3__0[22:22], termf_2[23:23], termf_1[23:23]);
  C3 I549 (fa3_23min_0[7:7], ct3__0[22:22], termf_2[23:23], termt_1[23:23]);
  NOR3 I550 (simp4151_0[0:0], fa3_23min_0[0:0], fa3_23min_0[3:3], fa3_23min_0[5:5]);
  INV I551 (simp4151_0[1:1], fa3_23min_0[6:6]);
  NAND2 I552 (o_0r0[23:23], simp4151_0[0:0], simp4151_0[1:1]);
  NOR3 I553 (simp4161_0[0:0], fa3_23min_0[1:1], fa3_23min_0[2:2], fa3_23min_0[4:4]);
  INV I554 (simp4161_0[1:1], fa3_23min_0[7:7]);
  NAND2 I555 (o_0r1[23:23], simp4161_0[0:0], simp4161_0[1:1]);
  AO222 I556 (ct3__0[23:23], termt_1[23:23], termf_2[23:23], termt_1[23:23], ct3__0[22:22], termf_2[23:23], ct3__0[22:22]);
  AO222 I557 (cf3__0[23:23], termf_1[23:23], termt_2[23:23], termf_1[23:23], cf3__0[22:22], termt_2[23:23], cf3__0[22:22]);
  C3 I558 (fa3_24min_0[0:0], cf3__0[23:23], termt_2[24:24], termf_1[24:24]);
  C3 I559 (fa3_24min_0[1:1], cf3__0[23:23], termt_2[24:24], termt_1[24:24]);
  C3 I560 (fa3_24min_0[2:2], cf3__0[23:23], termf_2[24:24], termf_1[24:24]);
  C3 I561 (fa3_24min_0[3:3], cf3__0[23:23], termf_2[24:24], termt_1[24:24]);
  C3 I562 (fa3_24min_0[4:4], ct3__0[23:23], termt_2[24:24], termf_1[24:24]);
  C3 I563 (fa3_24min_0[5:5], ct3__0[23:23], termt_2[24:24], termt_1[24:24]);
  C3 I564 (fa3_24min_0[6:6], ct3__0[23:23], termf_2[24:24], termf_1[24:24]);
  C3 I565 (fa3_24min_0[7:7], ct3__0[23:23], termf_2[24:24], termt_1[24:24]);
  NOR3 I566 (simp4281_0[0:0], fa3_24min_0[0:0], fa3_24min_0[3:3], fa3_24min_0[5:5]);
  INV I567 (simp4281_0[1:1], fa3_24min_0[6:6]);
  NAND2 I568 (o_0r0[24:24], simp4281_0[0:0], simp4281_0[1:1]);
  NOR3 I569 (simp4291_0[0:0], fa3_24min_0[1:1], fa3_24min_0[2:2], fa3_24min_0[4:4]);
  INV I570 (simp4291_0[1:1], fa3_24min_0[7:7]);
  NAND2 I571 (o_0r1[24:24], simp4291_0[0:0], simp4291_0[1:1]);
  AO222 I572 (ct3__0[24:24], termt_1[24:24], termf_2[24:24], termt_1[24:24], ct3__0[23:23], termf_2[24:24], ct3__0[23:23]);
  AO222 I573 (cf3__0[24:24], termf_1[24:24], termt_2[24:24], termf_1[24:24], cf3__0[23:23], termt_2[24:24], cf3__0[23:23]);
  C3 I574 (fa3_25min_0[0:0], cf3__0[24:24], termt_2[25:25], termf_1[25:25]);
  C3 I575 (fa3_25min_0[1:1], cf3__0[24:24], termt_2[25:25], termt_1[25:25]);
  C3 I576 (fa3_25min_0[2:2], cf3__0[24:24], termf_2[25:25], termf_1[25:25]);
  C3 I577 (fa3_25min_0[3:3], cf3__0[24:24], termf_2[25:25], termt_1[25:25]);
  C3 I578 (fa3_25min_0[4:4], ct3__0[24:24], termt_2[25:25], termf_1[25:25]);
  C3 I579 (fa3_25min_0[5:5], ct3__0[24:24], termt_2[25:25], termt_1[25:25]);
  C3 I580 (fa3_25min_0[6:6], ct3__0[24:24], termf_2[25:25], termf_1[25:25]);
  C3 I581 (fa3_25min_0[7:7], ct3__0[24:24], termf_2[25:25], termt_1[25:25]);
  NOR3 I582 (simp4411_0[0:0], fa3_25min_0[0:0], fa3_25min_0[3:3], fa3_25min_0[5:5]);
  INV I583 (simp4411_0[1:1], fa3_25min_0[6:6]);
  NAND2 I584 (o_0r0[25:25], simp4411_0[0:0], simp4411_0[1:1]);
  NOR3 I585 (simp4421_0[0:0], fa3_25min_0[1:1], fa3_25min_0[2:2], fa3_25min_0[4:4]);
  INV I586 (simp4421_0[1:1], fa3_25min_0[7:7]);
  NAND2 I587 (o_0r1[25:25], simp4421_0[0:0], simp4421_0[1:1]);
  AO222 I588 (ct3__0[25:25], termt_1[25:25], termf_2[25:25], termt_1[25:25], ct3__0[24:24], termf_2[25:25], ct3__0[24:24]);
  AO222 I589 (cf3__0[25:25], termf_1[25:25], termt_2[25:25], termf_1[25:25], cf3__0[24:24], termt_2[25:25], cf3__0[24:24]);
  C3 I590 (fa3_26min_0[0:0], cf3__0[25:25], termt_2[26:26], termf_1[26:26]);
  C3 I591 (fa3_26min_0[1:1], cf3__0[25:25], termt_2[26:26], termt_1[26:26]);
  C3 I592 (fa3_26min_0[2:2], cf3__0[25:25], termf_2[26:26], termf_1[26:26]);
  C3 I593 (fa3_26min_0[3:3], cf3__0[25:25], termf_2[26:26], termt_1[26:26]);
  C3 I594 (fa3_26min_0[4:4], ct3__0[25:25], termt_2[26:26], termf_1[26:26]);
  C3 I595 (fa3_26min_0[5:5], ct3__0[25:25], termt_2[26:26], termt_1[26:26]);
  C3 I596 (fa3_26min_0[6:6], ct3__0[25:25], termf_2[26:26], termf_1[26:26]);
  C3 I597 (fa3_26min_0[7:7], ct3__0[25:25], termf_2[26:26], termt_1[26:26]);
  NOR3 I598 (simp4541_0[0:0], fa3_26min_0[0:0], fa3_26min_0[3:3], fa3_26min_0[5:5]);
  INV I599 (simp4541_0[1:1], fa3_26min_0[6:6]);
  NAND2 I600 (o_0r0[26:26], simp4541_0[0:0], simp4541_0[1:1]);
  NOR3 I601 (simp4551_0[0:0], fa3_26min_0[1:1], fa3_26min_0[2:2], fa3_26min_0[4:4]);
  INV I602 (simp4551_0[1:1], fa3_26min_0[7:7]);
  NAND2 I603 (o_0r1[26:26], simp4551_0[0:0], simp4551_0[1:1]);
  AO222 I604 (ct3__0[26:26], termt_1[26:26], termf_2[26:26], termt_1[26:26], ct3__0[25:25], termf_2[26:26], ct3__0[25:25]);
  AO222 I605 (cf3__0[26:26], termf_1[26:26], termt_2[26:26], termf_1[26:26], cf3__0[25:25], termt_2[26:26], cf3__0[25:25]);
  C3 I606 (fa3_27min_0[0:0], cf3__0[26:26], termt_2[27:27], termf_1[27:27]);
  C3 I607 (fa3_27min_0[1:1], cf3__0[26:26], termt_2[27:27], termt_1[27:27]);
  C3 I608 (fa3_27min_0[2:2], cf3__0[26:26], termf_2[27:27], termf_1[27:27]);
  C3 I609 (fa3_27min_0[3:3], cf3__0[26:26], termf_2[27:27], termt_1[27:27]);
  C3 I610 (fa3_27min_0[4:4], ct3__0[26:26], termt_2[27:27], termf_1[27:27]);
  C3 I611 (fa3_27min_0[5:5], ct3__0[26:26], termt_2[27:27], termt_1[27:27]);
  C3 I612 (fa3_27min_0[6:6], ct3__0[26:26], termf_2[27:27], termf_1[27:27]);
  C3 I613 (fa3_27min_0[7:7], ct3__0[26:26], termf_2[27:27], termt_1[27:27]);
  NOR3 I614 (simp4671_0[0:0], fa3_27min_0[0:0], fa3_27min_0[3:3], fa3_27min_0[5:5]);
  INV I615 (simp4671_0[1:1], fa3_27min_0[6:6]);
  NAND2 I616 (o_0r0[27:27], simp4671_0[0:0], simp4671_0[1:1]);
  NOR3 I617 (simp4681_0[0:0], fa3_27min_0[1:1], fa3_27min_0[2:2], fa3_27min_0[4:4]);
  INV I618 (simp4681_0[1:1], fa3_27min_0[7:7]);
  NAND2 I619 (o_0r1[27:27], simp4681_0[0:0], simp4681_0[1:1]);
  AO222 I620 (ct3__0[27:27], termt_1[27:27], termf_2[27:27], termt_1[27:27], ct3__0[26:26], termf_2[27:27], ct3__0[26:26]);
  AO222 I621 (cf3__0[27:27], termf_1[27:27], termt_2[27:27], termf_1[27:27], cf3__0[26:26], termt_2[27:27], cf3__0[26:26]);
  C3 I622 (fa3_28min_0[0:0], cf3__0[27:27], termt_2[28:28], termf_1[28:28]);
  C3 I623 (fa3_28min_0[1:1], cf3__0[27:27], termt_2[28:28], termt_1[28:28]);
  C3 I624 (fa3_28min_0[2:2], cf3__0[27:27], termf_2[28:28], termf_1[28:28]);
  C3 I625 (fa3_28min_0[3:3], cf3__0[27:27], termf_2[28:28], termt_1[28:28]);
  C3 I626 (fa3_28min_0[4:4], ct3__0[27:27], termt_2[28:28], termf_1[28:28]);
  C3 I627 (fa3_28min_0[5:5], ct3__0[27:27], termt_2[28:28], termt_1[28:28]);
  C3 I628 (fa3_28min_0[6:6], ct3__0[27:27], termf_2[28:28], termf_1[28:28]);
  C3 I629 (fa3_28min_0[7:7], ct3__0[27:27], termf_2[28:28], termt_1[28:28]);
  NOR3 I630 (simp4801_0[0:0], fa3_28min_0[0:0], fa3_28min_0[3:3], fa3_28min_0[5:5]);
  INV I631 (simp4801_0[1:1], fa3_28min_0[6:6]);
  NAND2 I632 (o_0r0[28:28], simp4801_0[0:0], simp4801_0[1:1]);
  NOR3 I633 (simp4811_0[0:0], fa3_28min_0[1:1], fa3_28min_0[2:2], fa3_28min_0[4:4]);
  INV I634 (simp4811_0[1:1], fa3_28min_0[7:7]);
  NAND2 I635 (o_0r1[28:28], simp4811_0[0:0], simp4811_0[1:1]);
  AO222 I636 (ct3__0[28:28], termt_1[28:28], termf_2[28:28], termt_1[28:28], ct3__0[27:27], termf_2[28:28], ct3__0[27:27]);
  AO222 I637 (cf3__0[28:28], termf_1[28:28], termt_2[28:28], termf_1[28:28], cf3__0[27:27], termt_2[28:28], cf3__0[27:27]);
  C3 I638 (fa3_29min_0[0:0], cf3__0[28:28], termt_2[29:29], termf_1[29:29]);
  C3 I639 (fa3_29min_0[1:1], cf3__0[28:28], termt_2[29:29], termt_1[29:29]);
  C3 I640 (fa3_29min_0[2:2], cf3__0[28:28], termf_2[29:29], termf_1[29:29]);
  C3 I641 (fa3_29min_0[3:3], cf3__0[28:28], termf_2[29:29], termt_1[29:29]);
  C3 I642 (fa3_29min_0[4:4], ct3__0[28:28], termt_2[29:29], termf_1[29:29]);
  C3 I643 (fa3_29min_0[5:5], ct3__0[28:28], termt_2[29:29], termt_1[29:29]);
  C3 I644 (fa3_29min_0[6:6], ct3__0[28:28], termf_2[29:29], termf_1[29:29]);
  C3 I645 (fa3_29min_0[7:7], ct3__0[28:28], termf_2[29:29], termt_1[29:29]);
  NOR3 I646 (simp4931_0[0:0], fa3_29min_0[0:0], fa3_29min_0[3:3], fa3_29min_0[5:5]);
  INV I647 (simp4931_0[1:1], fa3_29min_0[6:6]);
  NAND2 I648 (o_0r0[29:29], simp4931_0[0:0], simp4931_0[1:1]);
  NOR3 I649 (simp4941_0[0:0], fa3_29min_0[1:1], fa3_29min_0[2:2], fa3_29min_0[4:4]);
  INV I650 (simp4941_0[1:1], fa3_29min_0[7:7]);
  NAND2 I651 (o_0r1[29:29], simp4941_0[0:0], simp4941_0[1:1]);
  AO222 I652 (ct3__0[29:29], termt_1[29:29], termf_2[29:29], termt_1[29:29], ct3__0[28:28], termf_2[29:29], ct3__0[28:28]);
  AO222 I653 (cf3__0[29:29], termf_1[29:29], termt_2[29:29], termf_1[29:29], cf3__0[28:28], termt_2[29:29], cf3__0[28:28]);
  C3 I654 (fa3_30min_0[0:0], cf3__0[29:29], termt_2[30:30], termf_1[30:30]);
  C3 I655 (fa3_30min_0[1:1], cf3__0[29:29], termt_2[30:30], termt_1[30:30]);
  C3 I656 (fa3_30min_0[2:2], cf3__0[29:29], termf_2[30:30], termf_1[30:30]);
  C3 I657 (fa3_30min_0[3:3], cf3__0[29:29], termf_2[30:30], termt_1[30:30]);
  C3 I658 (fa3_30min_0[4:4], ct3__0[29:29], termt_2[30:30], termf_1[30:30]);
  C3 I659 (fa3_30min_0[5:5], ct3__0[29:29], termt_2[30:30], termt_1[30:30]);
  C3 I660 (fa3_30min_0[6:6], ct3__0[29:29], termf_2[30:30], termf_1[30:30]);
  C3 I661 (fa3_30min_0[7:7], ct3__0[29:29], termf_2[30:30], termt_1[30:30]);
  NOR3 I662 (simp5061_0[0:0], fa3_30min_0[0:0], fa3_30min_0[3:3], fa3_30min_0[5:5]);
  INV I663 (simp5061_0[1:1], fa3_30min_0[6:6]);
  NAND2 I664 (o_0r0[30:30], simp5061_0[0:0], simp5061_0[1:1]);
  NOR3 I665 (simp5071_0[0:0], fa3_30min_0[1:1], fa3_30min_0[2:2], fa3_30min_0[4:4]);
  INV I666 (simp5071_0[1:1], fa3_30min_0[7:7]);
  NAND2 I667 (o_0r1[30:30], simp5071_0[0:0], simp5071_0[1:1]);
  AO222 I668 (ct3__0[30:30], termt_1[30:30], termf_2[30:30], termt_1[30:30], ct3__0[29:29], termf_2[30:30], ct3__0[29:29]);
  AO222 I669 (cf3__0[30:30], termf_1[30:30], termt_2[30:30], termf_1[30:30], cf3__0[29:29], termt_2[30:30], cf3__0[29:29]);
  C3 I670 (fa3_31min_0[0:0], cf3__0[30:30], termt_2[31:31], termf_1[31:31]);
  C3 I671 (fa3_31min_0[1:1], cf3__0[30:30], termt_2[31:31], termt_1[31:31]);
  C3 I672 (fa3_31min_0[2:2], cf3__0[30:30], termf_2[31:31], termf_1[31:31]);
  C3 I673 (fa3_31min_0[3:3], cf3__0[30:30], termf_2[31:31], termt_1[31:31]);
  C3 I674 (fa3_31min_0[4:4], ct3__0[30:30], termt_2[31:31], termf_1[31:31]);
  C3 I675 (fa3_31min_0[5:5], ct3__0[30:30], termt_2[31:31], termt_1[31:31]);
  C3 I676 (fa3_31min_0[6:6], ct3__0[30:30], termf_2[31:31], termf_1[31:31]);
  C3 I677 (fa3_31min_0[7:7], ct3__0[30:30], termf_2[31:31], termt_1[31:31]);
  NOR3 I678 (simp5191_0[0:0], fa3_31min_0[0:0], fa3_31min_0[3:3], fa3_31min_0[5:5]);
  INV I679 (simp5191_0[1:1], fa3_31min_0[6:6]);
  NAND2 I680 (o_0r0[31:31], simp5191_0[0:0], simp5191_0[1:1]);
  NOR3 I681 (simp5201_0[0:0], fa3_31min_0[1:1], fa3_31min_0[2:2], fa3_31min_0[4:4]);
  INV I682 (simp5201_0[1:1], fa3_31min_0[7:7]);
  NAND2 I683 (o_0r1[31:31], simp5201_0[0:0], simp5201_0[1:1]);
  AO222 I684 (ct3__0[31:31], termt_1[31:31], termf_2[31:31], termt_1[31:31], ct3__0[30:30], termf_2[31:31], ct3__0[30:30]);
  AO222 I685 (cf3__0[31:31], termf_1[31:31], termt_2[31:31], termf_1[31:31], cf3__0[30:30], termt_2[31:31], cf3__0[30:30]);
  C3 I686 (fa3_32min_0[0:0], cf3__0[31:31], termt_2[32:32], termf_1[32:32]);
  C3 I687 (fa3_32min_0[1:1], cf3__0[31:31], termt_2[32:32], termt_1[32:32]);
  C3 I688 (fa3_32min_0[2:2], cf3__0[31:31], termf_2[32:32], termf_1[32:32]);
  C3 I689 (fa3_32min_0[3:3], cf3__0[31:31], termf_2[32:32], termt_1[32:32]);
  C3 I690 (fa3_32min_0[4:4], ct3__0[31:31], termt_2[32:32], termf_1[32:32]);
  C3 I691 (fa3_32min_0[5:5], ct3__0[31:31], termt_2[32:32], termt_1[32:32]);
  C3 I692 (fa3_32min_0[6:6], ct3__0[31:31], termf_2[32:32], termf_1[32:32]);
  C3 I693 (fa3_32min_0[7:7], ct3__0[31:31], termf_2[32:32], termt_1[32:32]);
  NOR3 I694 (simp5321_0[0:0], fa3_32min_0[0:0], fa3_32min_0[3:3], fa3_32min_0[5:5]);
  INV I695 (simp5321_0[1:1], fa3_32min_0[6:6]);
  NAND2 I696 (o_0r0[32:32], simp5321_0[0:0], simp5321_0[1:1]);
  NOR3 I697 (simp5331_0[0:0], fa3_32min_0[1:1], fa3_32min_0[2:2], fa3_32min_0[4:4]);
  INV I698 (simp5331_0[1:1], fa3_32min_0[7:7]);
  NAND2 I699 (o_0r1[32:32], simp5331_0[0:0], simp5331_0[1:1]);
  AO222 I700 (ct3__0[32:32], termt_1[32:32], termf_2[32:32], termt_1[32:32], ct3__0[31:31], termf_2[32:32], ct3__0[31:31]);
  AO222 I701 (cf3__0[32:32], termf_1[32:32], termt_2[32:32], termf_1[32:32], cf3__0[31:31], termt_2[32:32], cf3__0[31:31]);
  BUFF I702 (i_0a, o_0a);
endmodule

// tko3m1_1nm3b1_2eqi0w3bt1o0w3b TeakO [
//     (1,TeakOConstant 3 1),
//     (2,TeakOp TeakOpEqual [(0,0+:3),(1,0+:3)])] [One 3,One 1]
module tko3m1_1nm3b1_2eqi0w3bt1o0w3b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [2:0] gocomp_0;
  wire [2:0] termf_1;
  wire [2:0] termt_1;
  wire [2:0] xf2_0;
  wire [2:0] xt2_0;
  wire [3:0] op2_0_0;
  wire [3:0] op2_1_0;
  wire [3:0] op2_2_0;
  wire [1:0] c2o_0;
  wire [1:0] c2o_1;
  wire [3:0] c2r0_0;
  wire [3:0] c20_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I3 (go_0, gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  BUFF I4 (termt_1[0:0], go_0);
  GND I5 (termf_1[0:0]);
  BUFF I6 (termf_1[1:1], go_0);
  BUFF I7 (termf_1[2:2], go_0);
  GND I8 (termt_1[1:1]);
  GND I9 (termt_1[2:2]);
  C2 I10 (op2_0_0[0:0], termf_1[0:0], i_0r0[0:0]);
  C2 I11 (op2_0_0[1:1], termf_1[0:0], i_0r1[0:0]);
  C2 I12 (op2_0_0[2:2], termt_1[0:0], i_0r0[0:0]);
  C2 I13 (op2_0_0[3:3], termt_1[0:0], i_0r1[0:0]);
  OR2 I14 (xf2_0[0:0], op2_0_0[1:1], op2_0_0[2:2]);
  OR2 I15 (xt2_0[0:0], op2_0_0[0:0], op2_0_0[3:3]);
  C2 I16 (op2_1_0[0:0], termf_1[1:1], i_0r0[1:1]);
  C2 I17 (op2_1_0[1:1], termf_1[1:1], i_0r1[1:1]);
  C2 I18 (op2_1_0[2:2], termt_1[1:1], i_0r0[1:1]);
  C2 I19 (op2_1_0[3:3], termt_1[1:1], i_0r1[1:1]);
  OR2 I20 (xf2_0[1:1], op2_1_0[1:1], op2_1_0[2:2]);
  OR2 I21 (xt2_0[1:1], op2_1_0[0:0], op2_1_0[3:3]);
  C2 I22 (op2_2_0[0:0], termf_1[2:2], i_0r0[2:2]);
  C2 I23 (op2_2_0[1:1], termf_1[2:2], i_0r1[2:2]);
  C2 I24 (op2_2_0[2:2], termt_1[2:2], i_0r0[2:2]);
  C2 I25 (op2_2_0[3:3], termt_1[2:2], i_0r1[2:2]);
  OR2 I26 (xf2_0[2:2], op2_2_0[1:1], op2_2_0[2:2]);
  OR2 I27 (xt2_0[2:2], op2_2_0[0:0], op2_2_0[3:3]);
  C2 I28 (c2r0_0[0:0], c2o_0[1:1], c2o_0[0:0]);
  C2 I29 (c2r0_0[1:1], c2o_0[1:1], c2o_1[0:0]);
  C2 I30 (c2r0_0[2:2], c2o_1[1:1], c2o_0[0:0]);
  C2 I31 (c2r0_0[3:3], c2o_1[1:1], c2o_1[0:0]);
  OR3 I32 (o_0r0, c2r0_0[0:0], c2r0_0[1:1], c2r0_0[2:2]);
  BUFF I33 (o_0r1, c2r0_0[3:3]);
  BUFF I34 (c2o_0[1:1], xf2_0[2:2]);
  BUFF I35 (c2o_1[1:1], xt2_0[2:2]);
  C2 I36 (c20_0[0:0], xf2_0[1:1], xf2_0[0:0]);
  C2 I37 (c20_0[1:1], xf2_0[1:1], xt2_0[0:0]);
  C2 I38 (c20_0[2:2], xt2_0[1:1], xf2_0[0:0]);
  C2 I39 (c20_0[3:3], xt2_0[1:1], xt2_0[0:0]);
  OR3 I40 (c2o_0[0:0], c20_0[0:0], c20_0[1:1], c20_0[2:2]);
  BUFF I41 (c2o_1[0:0], c20_0[3:3]);
  BUFF I42 (i_0a, o_0a);
endmodule

// tkj32m32_0_0_0 TeakJ [Many [32,0,0,0],One 32]
module tkj32m32_0_0_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_0r1[24:24]);
  BUFF I57 (joint_0[25:25], i_0r1[25:25]);
  BUFF I58 (joint_0[26:26], i_0r1[26:26]);
  BUFF I59 (joint_0[27:27], i_0r1[27:27]);
  BUFF I60 (joint_0[28:28], i_0r1[28:28]);
  BUFF I61 (joint_0[29:29], i_0r1[29:29]);
  BUFF I62 (joint_0[30:30], i_0r1[30:30]);
  BUFF I63 (joint_0[31:31], i_0r1[31:31]);
  C3 I64 (icomplete_0, i_1r, i_2r, i_3r);
  C2 I65 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I66 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I67 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I68 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I69 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I70 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I71 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I72 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I73 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I74 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I75 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I76 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I77 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I78 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I79 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I80 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I81 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I82 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I83 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I84 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I85 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I86 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I87 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I88 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I89 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I90 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I91 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I92 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I93 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I94 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I95 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I96 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I97 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I98 (o_0r1[1:1], joint_0[1:1]);
  BUFF I99 (o_0r1[2:2], joint_0[2:2]);
  BUFF I100 (o_0r1[3:3], joint_0[3:3]);
  BUFF I101 (o_0r1[4:4], joint_0[4:4]);
  BUFF I102 (o_0r1[5:5], joint_0[5:5]);
  BUFF I103 (o_0r1[6:6], joint_0[6:6]);
  BUFF I104 (o_0r1[7:7], joint_0[7:7]);
  BUFF I105 (o_0r1[8:8], joint_0[8:8]);
  BUFF I106 (o_0r1[9:9], joint_0[9:9]);
  BUFF I107 (o_0r1[10:10], joint_0[10:10]);
  BUFF I108 (o_0r1[11:11], joint_0[11:11]);
  BUFF I109 (o_0r1[12:12], joint_0[12:12]);
  BUFF I110 (o_0r1[13:13], joint_0[13:13]);
  BUFF I111 (o_0r1[14:14], joint_0[14:14]);
  BUFF I112 (o_0r1[15:15], joint_0[15:15]);
  BUFF I113 (o_0r1[16:16], joint_0[16:16]);
  BUFF I114 (o_0r1[17:17], joint_0[17:17]);
  BUFF I115 (o_0r1[18:18], joint_0[18:18]);
  BUFF I116 (o_0r1[19:19], joint_0[19:19]);
  BUFF I117 (o_0r1[20:20], joint_0[20:20]);
  BUFF I118 (o_0r1[21:21], joint_0[21:21]);
  BUFF I119 (o_0r1[22:22], joint_0[22:22]);
  BUFF I120 (o_0r1[23:23], joint_0[23:23]);
  BUFF I121 (o_0r1[24:24], joint_0[24:24]);
  BUFF I122 (o_0r1[25:25], joint_0[25:25]);
  BUFF I123 (o_0r1[26:26], joint_0[26:26]);
  BUFF I124 (o_0r1[27:27], joint_0[27:27]);
  BUFF I125 (o_0r1[28:28], joint_0[28:28]);
  BUFF I126 (o_0r1[29:29], joint_0[29:29]);
  BUFF I127 (o_0r1[30:30], joint_0[30:30]);
  BUFF I128 (o_0r1[31:31], joint_0[31:31]);
  BUFF I129 (i_0a, o_0a);
  BUFF I130 (i_1a, o_0a);
  BUFF I131 (i_2a, o_0a);
  BUFF I132 (i_3a, o_0a);
endmodule

// tko64m32_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b_4apt3o0w32b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32),(0,31+:1)]),
//     (2,TeakOAppend 1 [(0,32+:32),(0,63+:1)]),
//     (3,TeakOp TeakOpAdd [(1,0+:33),(2,0+:33)]),
//     (4,TeakOAppend 1 [(3,0+:32)])] [One 64,One 32]
module tko64m32_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b_4apt3o0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [32:0] termf_1;
  wire [32:0] termf_2;
  wire [32:0] termf_3;
  wire [32:0] termt_1;
  wire [32:0] termt_2;
  wire [32:0] termt_3;
  wire [32:0] cf3__0;
  wire [32:0] ct3__0;
  wire [3:0] ha3__0;
  wire [7:0] fa3_1min_0;
  wire [1:0] simp1581_0;
  wire [1:0] simp1591_0;
  wire [7:0] fa3_2min_0;
  wire [1:0] simp1711_0;
  wire [1:0] simp1721_0;
  wire [7:0] fa3_3min_0;
  wire [1:0] simp1841_0;
  wire [1:0] simp1851_0;
  wire [7:0] fa3_4min_0;
  wire [1:0] simp1971_0;
  wire [1:0] simp1981_0;
  wire [7:0] fa3_5min_0;
  wire [1:0] simp2101_0;
  wire [1:0] simp2111_0;
  wire [7:0] fa3_6min_0;
  wire [1:0] simp2231_0;
  wire [1:0] simp2241_0;
  wire [7:0] fa3_7min_0;
  wire [1:0] simp2361_0;
  wire [1:0] simp2371_0;
  wire [7:0] fa3_8min_0;
  wire [1:0] simp2491_0;
  wire [1:0] simp2501_0;
  wire [7:0] fa3_9min_0;
  wire [1:0] simp2621_0;
  wire [1:0] simp2631_0;
  wire [7:0] fa3_10min_0;
  wire [1:0] simp2751_0;
  wire [1:0] simp2761_0;
  wire [7:0] fa3_11min_0;
  wire [1:0] simp2881_0;
  wire [1:0] simp2891_0;
  wire [7:0] fa3_12min_0;
  wire [1:0] simp3011_0;
  wire [1:0] simp3021_0;
  wire [7:0] fa3_13min_0;
  wire [1:0] simp3141_0;
  wire [1:0] simp3151_0;
  wire [7:0] fa3_14min_0;
  wire [1:0] simp3271_0;
  wire [1:0] simp3281_0;
  wire [7:0] fa3_15min_0;
  wire [1:0] simp3401_0;
  wire [1:0] simp3411_0;
  wire [7:0] fa3_16min_0;
  wire [1:0] simp3531_0;
  wire [1:0] simp3541_0;
  wire [7:0] fa3_17min_0;
  wire [1:0] simp3661_0;
  wire [1:0] simp3671_0;
  wire [7:0] fa3_18min_0;
  wire [1:0] simp3791_0;
  wire [1:0] simp3801_0;
  wire [7:0] fa3_19min_0;
  wire [1:0] simp3921_0;
  wire [1:0] simp3931_0;
  wire [7:0] fa3_20min_0;
  wire [1:0] simp4051_0;
  wire [1:0] simp4061_0;
  wire [7:0] fa3_21min_0;
  wire [1:0] simp4181_0;
  wire [1:0] simp4191_0;
  wire [7:0] fa3_22min_0;
  wire [1:0] simp4311_0;
  wire [1:0] simp4321_0;
  wire [7:0] fa3_23min_0;
  wire [1:0] simp4441_0;
  wire [1:0] simp4451_0;
  wire [7:0] fa3_24min_0;
  wire [1:0] simp4571_0;
  wire [1:0] simp4581_0;
  wire [7:0] fa3_25min_0;
  wire [1:0] simp4701_0;
  wire [1:0] simp4711_0;
  wire [7:0] fa3_26min_0;
  wire [1:0] simp4831_0;
  wire [1:0] simp4841_0;
  wire [7:0] fa3_27min_0;
  wire [1:0] simp4961_0;
  wire [1:0] simp4971_0;
  wire [7:0] fa3_28min_0;
  wire [1:0] simp5091_0;
  wire [1:0] simp5101_0;
  wire [7:0] fa3_29min_0;
  wire [1:0] simp5221_0;
  wire [1:0] simp5231_0;
  wire [7:0] fa3_30min_0;
  wire [1:0] simp5351_0;
  wire [1:0] simp5361_0;
  wire [7:0] fa3_31min_0;
  wire [1:0] simp5481_0;
  wire [1:0] simp5491_0;
  wire [7:0] fa3_32min_0;
  wire [1:0] simp5611_0;
  wire [1:0] simp5621_0;
  BUFF I0 (termf_1[0:0], i_0r0[0:0]);
  BUFF I1 (termf_1[1:1], i_0r0[1:1]);
  BUFF I2 (termf_1[2:2], i_0r0[2:2]);
  BUFF I3 (termf_1[3:3], i_0r0[3:3]);
  BUFF I4 (termf_1[4:4], i_0r0[4:4]);
  BUFF I5 (termf_1[5:5], i_0r0[5:5]);
  BUFF I6 (termf_1[6:6], i_0r0[6:6]);
  BUFF I7 (termf_1[7:7], i_0r0[7:7]);
  BUFF I8 (termf_1[8:8], i_0r0[8:8]);
  BUFF I9 (termf_1[9:9], i_0r0[9:9]);
  BUFF I10 (termf_1[10:10], i_0r0[10:10]);
  BUFF I11 (termf_1[11:11], i_0r0[11:11]);
  BUFF I12 (termf_1[12:12], i_0r0[12:12]);
  BUFF I13 (termf_1[13:13], i_0r0[13:13]);
  BUFF I14 (termf_1[14:14], i_0r0[14:14]);
  BUFF I15 (termf_1[15:15], i_0r0[15:15]);
  BUFF I16 (termf_1[16:16], i_0r0[16:16]);
  BUFF I17 (termf_1[17:17], i_0r0[17:17]);
  BUFF I18 (termf_1[18:18], i_0r0[18:18]);
  BUFF I19 (termf_1[19:19], i_0r0[19:19]);
  BUFF I20 (termf_1[20:20], i_0r0[20:20]);
  BUFF I21 (termf_1[21:21], i_0r0[21:21]);
  BUFF I22 (termf_1[22:22], i_0r0[22:22]);
  BUFF I23 (termf_1[23:23], i_0r0[23:23]);
  BUFF I24 (termf_1[24:24], i_0r0[24:24]);
  BUFF I25 (termf_1[25:25], i_0r0[25:25]);
  BUFF I26 (termf_1[26:26], i_0r0[26:26]);
  BUFF I27 (termf_1[27:27], i_0r0[27:27]);
  BUFF I28 (termf_1[28:28], i_0r0[28:28]);
  BUFF I29 (termf_1[29:29], i_0r0[29:29]);
  BUFF I30 (termf_1[30:30], i_0r0[30:30]);
  BUFF I31 (termf_1[31:31], i_0r0[31:31]);
  BUFF I32 (termf_1[32:32], i_0r0[31:31]);
  BUFF I33 (termt_1[0:0], i_0r1[0:0]);
  BUFF I34 (termt_1[1:1], i_0r1[1:1]);
  BUFF I35 (termt_1[2:2], i_0r1[2:2]);
  BUFF I36 (termt_1[3:3], i_0r1[3:3]);
  BUFF I37 (termt_1[4:4], i_0r1[4:4]);
  BUFF I38 (termt_1[5:5], i_0r1[5:5]);
  BUFF I39 (termt_1[6:6], i_0r1[6:6]);
  BUFF I40 (termt_1[7:7], i_0r1[7:7]);
  BUFF I41 (termt_1[8:8], i_0r1[8:8]);
  BUFF I42 (termt_1[9:9], i_0r1[9:9]);
  BUFF I43 (termt_1[10:10], i_0r1[10:10]);
  BUFF I44 (termt_1[11:11], i_0r1[11:11]);
  BUFF I45 (termt_1[12:12], i_0r1[12:12]);
  BUFF I46 (termt_1[13:13], i_0r1[13:13]);
  BUFF I47 (termt_1[14:14], i_0r1[14:14]);
  BUFF I48 (termt_1[15:15], i_0r1[15:15]);
  BUFF I49 (termt_1[16:16], i_0r1[16:16]);
  BUFF I50 (termt_1[17:17], i_0r1[17:17]);
  BUFF I51 (termt_1[18:18], i_0r1[18:18]);
  BUFF I52 (termt_1[19:19], i_0r1[19:19]);
  BUFF I53 (termt_1[20:20], i_0r1[20:20]);
  BUFF I54 (termt_1[21:21], i_0r1[21:21]);
  BUFF I55 (termt_1[22:22], i_0r1[22:22]);
  BUFF I56 (termt_1[23:23], i_0r1[23:23]);
  BUFF I57 (termt_1[24:24], i_0r1[24:24]);
  BUFF I58 (termt_1[25:25], i_0r1[25:25]);
  BUFF I59 (termt_1[26:26], i_0r1[26:26]);
  BUFF I60 (termt_1[27:27], i_0r1[27:27]);
  BUFF I61 (termt_1[28:28], i_0r1[28:28]);
  BUFF I62 (termt_1[29:29], i_0r1[29:29]);
  BUFF I63 (termt_1[30:30], i_0r1[30:30]);
  BUFF I64 (termt_1[31:31], i_0r1[31:31]);
  BUFF I65 (termt_1[32:32], i_0r1[31:31]);
  BUFF I66 (termf_2[0:0], i_0r0[32:32]);
  BUFF I67 (termf_2[1:1], i_0r0[33:33]);
  BUFF I68 (termf_2[2:2], i_0r0[34:34]);
  BUFF I69 (termf_2[3:3], i_0r0[35:35]);
  BUFF I70 (termf_2[4:4], i_0r0[36:36]);
  BUFF I71 (termf_2[5:5], i_0r0[37:37]);
  BUFF I72 (termf_2[6:6], i_0r0[38:38]);
  BUFF I73 (termf_2[7:7], i_0r0[39:39]);
  BUFF I74 (termf_2[8:8], i_0r0[40:40]);
  BUFF I75 (termf_2[9:9], i_0r0[41:41]);
  BUFF I76 (termf_2[10:10], i_0r0[42:42]);
  BUFF I77 (termf_2[11:11], i_0r0[43:43]);
  BUFF I78 (termf_2[12:12], i_0r0[44:44]);
  BUFF I79 (termf_2[13:13], i_0r0[45:45]);
  BUFF I80 (termf_2[14:14], i_0r0[46:46]);
  BUFF I81 (termf_2[15:15], i_0r0[47:47]);
  BUFF I82 (termf_2[16:16], i_0r0[48:48]);
  BUFF I83 (termf_2[17:17], i_0r0[49:49]);
  BUFF I84 (termf_2[18:18], i_0r0[50:50]);
  BUFF I85 (termf_2[19:19], i_0r0[51:51]);
  BUFF I86 (termf_2[20:20], i_0r0[52:52]);
  BUFF I87 (termf_2[21:21], i_0r0[53:53]);
  BUFF I88 (termf_2[22:22], i_0r0[54:54]);
  BUFF I89 (termf_2[23:23], i_0r0[55:55]);
  BUFF I90 (termf_2[24:24], i_0r0[56:56]);
  BUFF I91 (termf_2[25:25], i_0r0[57:57]);
  BUFF I92 (termf_2[26:26], i_0r0[58:58]);
  BUFF I93 (termf_2[27:27], i_0r0[59:59]);
  BUFF I94 (termf_2[28:28], i_0r0[60:60]);
  BUFF I95 (termf_2[29:29], i_0r0[61:61]);
  BUFF I96 (termf_2[30:30], i_0r0[62:62]);
  BUFF I97 (termf_2[31:31], i_0r0[63:63]);
  BUFF I98 (termf_2[32:32], i_0r0[63:63]);
  BUFF I99 (termt_2[0:0], i_0r1[32:32]);
  BUFF I100 (termt_2[1:1], i_0r1[33:33]);
  BUFF I101 (termt_2[2:2], i_0r1[34:34]);
  BUFF I102 (termt_2[3:3], i_0r1[35:35]);
  BUFF I103 (termt_2[4:4], i_0r1[36:36]);
  BUFF I104 (termt_2[5:5], i_0r1[37:37]);
  BUFF I105 (termt_2[6:6], i_0r1[38:38]);
  BUFF I106 (termt_2[7:7], i_0r1[39:39]);
  BUFF I107 (termt_2[8:8], i_0r1[40:40]);
  BUFF I108 (termt_2[9:9], i_0r1[41:41]);
  BUFF I109 (termt_2[10:10], i_0r1[42:42]);
  BUFF I110 (termt_2[11:11], i_0r1[43:43]);
  BUFF I111 (termt_2[12:12], i_0r1[44:44]);
  BUFF I112 (termt_2[13:13], i_0r1[45:45]);
  BUFF I113 (termt_2[14:14], i_0r1[46:46]);
  BUFF I114 (termt_2[15:15], i_0r1[47:47]);
  BUFF I115 (termt_2[16:16], i_0r1[48:48]);
  BUFF I116 (termt_2[17:17], i_0r1[49:49]);
  BUFF I117 (termt_2[18:18], i_0r1[50:50]);
  BUFF I118 (termt_2[19:19], i_0r1[51:51]);
  BUFF I119 (termt_2[20:20], i_0r1[52:52]);
  BUFF I120 (termt_2[21:21], i_0r1[53:53]);
  BUFF I121 (termt_2[22:22], i_0r1[54:54]);
  BUFF I122 (termt_2[23:23], i_0r1[55:55]);
  BUFF I123 (termt_2[24:24], i_0r1[56:56]);
  BUFF I124 (termt_2[25:25], i_0r1[57:57]);
  BUFF I125 (termt_2[26:26], i_0r1[58:58]);
  BUFF I126 (termt_2[27:27], i_0r1[59:59]);
  BUFF I127 (termt_2[28:28], i_0r1[60:60]);
  BUFF I128 (termt_2[29:29], i_0r1[61:61]);
  BUFF I129 (termt_2[30:30], i_0r1[62:62]);
  BUFF I130 (termt_2[31:31], i_0r1[63:63]);
  BUFF I131 (termt_2[32:32], i_0r1[63:63]);
  C2 I132 (ha3__0[0:0], termf_2[0:0], termf_1[0:0]);
  C2 I133 (ha3__0[1:1], termf_2[0:0], termt_1[0:0]);
  C2 I134 (ha3__0[2:2], termt_2[0:0], termf_1[0:0]);
  C2 I135 (ha3__0[3:3], termt_2[0:0], termt_1[0:0]);
  OR3 I136 (cf3__0[0:0], ha3__0[0:0], ha3__0[1:1], ha3__0[2:2]);
  BUFF I137 (ct3__0[0:0], ha3__0[3:3]);
  OR2 I138 (termf_3[0:0], ha3__0[0:0], ha3__0[3:3]);
  OR2 I139 (termt_3[0:0], ha3__0[1:1], ha3__0[2:2]);
  C3 I140 (fa3_1min_0[0:0], cf3__0[0:0], termf_2[1:1], termf_1[1:1]);
  C3 I141 (fa3_1min_0[1:1], cf3__0[0:0], termf_2[1:1], termt_1[1:1]);
  C3 I142 (fa3_1min_0[2:2], cf3__0[0:0], termt_2[1:1], termf_1[1:1]);
  C3 I143 (fa3_1min_0[3:3], cf3__0[0:0], termt_2[1:1], termt_1[1:1]);
  C3 I144 (fa3_1min_0[4:4], ct3__0[0:0], termf_2[1:1], termf_1[1:1]);
  C3 I145 (fa3_1min_0[5:5], ct3__0[0:0], termf_2[1:1], termt_1[1:1]);
  C3 I146 (fa3_1min_0[6:6], ct3__0[0:0], termt_2[1:1], termf_1[1:1]);
  C3 I147 (fa3_1min_0[7:7], ct3__0[0:0], termt_2[1:1], termt_1[1:1]);
  NOR3 I148 (simp1581_0[0:0], fa3_1min_0[0:0], fa3_1min_0[3:3], fa3_1min_0[5:5]);
  INV I149 (simp1581_0[1:1], fa3_1min_0[6:6]);
  NAND2 I150 (termf_3[1:1], simp1581_0[0:0], simp1581_0[1:1]);
  NOR3 I151 (simp1591_0[0:0], fa3_1min_0[1:1], fa3_1min_0[2:2], fa3_1min_0[4:4]);
  INV I152 (simp1591_0[1:1], fa3_1min_0[7:7]);
  NAND2 I153 (termt_3[1:1], simp1591_0[0:0], simp1591_0[1:1]);
  AO222 I154 (ct3__0[1:1], termt_1[1:1], termt_2[1:1], termt_1[1:1], ct3__0[0:0], termt_2[1:1], ct3__0[0:0]);
  AO222 I155 (cf3__0[1:1], termf_1[1:1], termf_2[1:1], termf_1[1:1], cf3__0[0:0], termf_2[1:1], cf3__0[0:0]);
  C3 I156 (fa3_2min_0[0:0], cf3__0[1:1], termf_2[2:2], termf_1[2:2]);
  C3 I157 (fa3_2min_0[1:1], cf3__0[1:1], termf_2[2:2], termt_1[2:2]);
  C3 I158 (fa3_2min_0[2:2], cf3__0[1:1], termt_2[2:2], termf_1[2:2]);
  C3 I159 (fa3_2min_0[3:3], cf3__0[1:1], termt_2[2:2], termt_1[2:2]);
  C3 I160 (fa3_2min_0[4:4], ct3__0[1:1], termf_2[2:2], termf_1[2:2]);
  C3 I161 (fa3_2min_0[5:5], ct3__0[1:1], termf_2[2:2], termt_1[2:2]);
  C3 I162 (fa3_2min_0[6:6], ct3__0[1:1], termt_2[2:2], termf_1[2:2]);
  C3 I163 (fa3_2min_0[7:7], ct3__0[1:1], termt_2[2:2], termt_1[2:2]);
  NOR3 I164 (simp1711_0[0:0], fa3_2min_0[0:0], fa3_2min_0[3:3], fa3_2min_0[5:5]);
  INV I165 (simp1711_0[1:1], fa3_2min_0[6:6]);
  NAND2 I166 (termf_3[2:2], simp1711_0[0:0], simp1711_0[1:1]);
  NOR3 I167 (simp1721_0[0:0], fa3_2min_0[1:1], fa3_2min_0[2:2], fa3_2min_0[4:4]);
  INV I168 (simp1721_0[1:1], fa3_2min_0[7:7]);
  NAND2 I169 (termt_3[2:2], simp1721_0[0:0], simp1721_0[1:1]);
  AO222 I170 (ct3__0[2:2], termt_1[2:2], termt_2[2:2], termt_1[2:2], ct3__0[1:1], termt_2[2:2], ct3__0[1:1]);
  AO222 I171 (cf3__0[2:2], termf_1[2:2], termf_2[2:2], termf_1[2:2], cf3__0[1:1], termf_2[2:2], cf3__0[1:1]);
  C3 I172 (fa3_3min_0[0:0], cf3__0[2:2], termf_2[3:3], termf_1[3:3]);
  C3 I173 (fa3_3min_0[1:1], cf3__0[2:2], termf_2[3:3], termt_1[3:3]);
  C3 I174 (fa3_3min_0[2:2], cf3__0[2:2], termt_2[3:3], termf_1[3:3]);
  C3 I175 (fa3_3min_0[3:3], cf3__0[2:2], termt_2[3:3], termt_1[3:3]);
  C3 I176 (fa3_3min_0[4:4], ct3__0[2:2], termf_2[3:3], termf_1[3:3]);
  C3 I177 (fa3_3min_0[5:5], ct3__0[2:2], termf_2[3:3], termt_1[3:3]);
  C3 I178 (fa3_3min_0[6:6], ct3__0[2:2], termt_2[3:3], termf_1[3:3]);
  C3 I179 (fa3_3min_0[7:7], ct3__0[2:2], termt_2[3:3], termt_1[3:3]);
  NOR3 I180 (simp1841_0[0:0], fa3_3min_0[0:0], fa3_3min_0[3:3], fa3_3min_0[5:5]);
  INV I181 (simp1841_0[1:1], fa3_3min_0[6:6]);
  NAND2 I182 (termf_3[3:3], simp1841_0[0:0], simp1841_0[1:1]);
  NOR3 I183 (simp1851_0[0:0], fa3_3min_0[1:1], fa3_3min_0[2:2], fa3_3min_0[4:4]);
  INV I184 (simp1851_0[1:1], fa3_3min_0[7:7]);
  NAND2 I185 (termt_3[3:3], simp1851_0[0:0], simp1851_0[1:1]);
  AO222 I186 (ct3__0[3:3], termt_1[3:3], termt_2[3:3], termt_1[3:3], ct3__0[2:2], termt_2[3:3], ct3__0[2:2]);
  AO222 I187 (cf3__0[3:3], termf_1[3:3], termf_2[3:3], termf_1[3:3], cf3__0[2:2], termf_2[3:3], cf3__0[2:2]);
  C3 I188 (fa3_4min_0[0:0], cf3__0[3:3], termf_2[4:4], termf_1[4:4]);
  C3 I189 (fa3_4min_0[1:1], cf3__0[3:3], termf_2[4:4], termt_1[4:4]);
  C3 I190 (fa3_4min_0[2:2], cf3__0[3:3], termt_2[4:4], termf_1[4:4]);
  C3 I191 (fa3_4min_0[3:3], cf3__0[3:3], termt_2[4:4], termt_1[4:4]);
  C3 I192 (fa3_4min_0[4:4], ct3__0[3:3], termf_2[4:4], termf_1[4:4]);
  C3 I193 (fa3_4min_0[5:5], ct3__0[3:3], termf_2[4:4], termt_1[4:4]);
  C3 I194 (fa3_4min_0[6:6], ct3__0[3:3], termt_2[4:4], termf_1[4:4]);
  C3 I195 (fa3_4min_0[7:7], ct3__0[3:3], termt_2[4:4], termt_1[4:4]);
  NOR3 I196 (simp1971_0[0:0], fa3_4min_0[0:0], fa3_4min_0[3:3], fa3_4min_0[5:5]);
  INV I197 (simp1971_0[1:1], fa3_4min_0[6:6]);
  NAND2 I198 (termf_3[4:4], simp1971_0[0:0], simp1971_0[1:1]);
  NOR3 I199 (simp1981_0[0:0], fa3_4min_0[1:1], fa3_4min_0[2:2], fa3_4min_0[4:4]);
  INV I200 (simp1981_0[1:1], fa3_4min_0[7:7]);
  NAND2 I201 (termt_3[4:4], simp1981_0[0:0], simp1981_0[1:1]);
  AO222 I202 (ct3__0[4:4], termt_1[4:4], termt_2[4:4], termt_1[4:4], ct3__0[3:3], termt_2[4:4], ct3__0[3:3]);
  AO222 I203 (cf3__0[4:4], termf_1[4:4], termf_2[4:4], termf_1[4:4], cf3__0[3:3], termf_2[4:4], cf3__0[3:3]);
  C3 I204 (fa3_5min_0[0:0], cf3__0[4:4], termf_2[5:5], termf_1[5:5]);
  C3 I205 (fa3_5min_0[1:1], cf3__0[4:4], termf_2[5:5], termt_1[5:5]);
  C3 I206 (fa3_5min_0[2:2], cf3__0[4:4], termt_2[5:5], termf_1[5:5]);
  C3 I207 (fa3_5min_0[3:3], cf3__0[4:4], termt_2[5:5], termt_1[5:5]);
  C3 I208 (fa3_5min_0[4:4], ct3__0[4:4], termf_2[5:5], termf_1[5:5]);
  C3 I209 (fa3_5min_0[5:5], ct3__0[4:4], termf_2[5:5], termt_1[5:5]);
  C3 I210 (fa3_5min_0[6:6], ct3__0[4:4], termt_2[5:5], termf_1[5:5]);
  C3 I211 (fa3_5min_0[7:7], ct3__0[4:4], termt_2[5:5], termt_1[5:5]);
  NOR3 I212 (simp2101_0[0:0], fa3_5min_0[0:0], fa3_5min_0[3:3], fa3_5min_0[5:5]);
  INV I213 (simp2101_0[1:1], fa3_5min_0[6:6]);
  NAND2 I214 (termf_3[5:5], simp2101_0[0:0], simp2101_0[1:1]);
  NOR3 I215 (simp2111_0[0:0], fa3_5min_0[1:1], fa3_5min_0[2:2], fa3_5min_0[4:4]);
  INV I216 (simp2111_0[1:1], fa3_5min_0[7:7]);
  NAND2 I217 (termt_3[5:5], simp2111_0[0:0], simp2111_0[1:1]);
  AO222 I218 (ct3__0[5:5], termt_1[5:5], termt_2[5:5], termt_1[5:5], ct3__0[4:4], termt_2[5:5], ct3__0[4:4]);
  AO222 I219 (cf3__0[5:5], termf_1[5:5], termf_2[5:5], termf_1[5:5], cf3__0[4:4], termf_2[5:5], cf3__0[4:4]);
  C3 I220 (fa3_6min_0[0:0], cf3__0[5:5], termf_2[6:6], termf_1[6:6]);
  C3 I221 (fa3_6min_0[1:1], cf3__0[5:5], termf_2[6:6], termt_1[6:6]);
  C3 I222 (fa3_6min_0[2:2], cf3__0[5:5], termt_2[6:6], termf_1[6:6]);
  C3 I223 (fa3_6min_0[3:3], cf3__0[5:5], termt_2[6:6], termt_1[6:6]);
  C3 I224 (fa3_6min_0[4:4], ct3__0[5:5], termf_2[6:6], termf_1[6:6]);
  C3 I225 (fa3_6min_0[5:5], ct3__0[5:5], termf_2[6:6], termt_1[6:6]);
  C3 I226 (fa3_6min_0[6:6], ct3__0[5:5], termt_2[6:6], termf_1[6:6]);
  C3 I227 (fa3_6min_0[7:7], ct3__0[5:5], termt_2[6:6], termt_1[6:6]);
  NOR3 I228 (simp2231_0[0:0], fa3_6min_0[0:0], fa3_6min_0[3:3], fa3_6min_0[5:5]);
  INV I229 (simp2231_0[1:1], fa3_6min_0[6:6]);
  NAND2 I230 (termf_3[6:6], simp2231_0[0:0], simp2231_0[1:1]);
  NOR3 I231 (simp2241_0[0:0], fa3_6min_0[1:1], fa3_6min_0[2:2], fa3_6min_0[4:4]);
  INV I232 (simp2241_0[1:1], fa3_6min_0[7:7]);
  NAND2 I233 (termt_3[6:6], simp2241_0[0:0], simp2241_0[1:1]);
  AO222 I234 (ct3__0[6:6], termt_1[6:6], termt_2[6:6], termt_1[6:6], ct3__0[5:5], termt_2[6:6], ct3__0[5:5]);
  AO222 I235 (cf3__0[6:6], termf_1[6:6], termf_2[6:6], termf_1[6:6], cf3__0[5:5], termf_2[6:6], cf3__0[5:5]);
  C3 I236 (fa3_7min_0[0:0], cf3__0[6:6], termf_2[7:7], termf_1[7:7]);
  C3 I237 (fa3_7min_0[1:1], cf3__0[6:6], termf_2[7:7], termt_1[7:7]);
  C3 I238 (fa3_7min_0[2:2], cf3__0[6:6], termt_2[7:7], termf_1[7:7]);
  C3 I239 (fa3_7min_0[3:3], cf3__0[6:6], termt_2[7:7], termt_1[7:7]);
  C3 I240 (fa3_7min_0[4:4], ct3__0[6:6], termf_2[7:7], termf_1[7:7]);
  C3 I241 (fa3_7min_0[5:5], ct3__0[6:6], termf_2[7:7], termt_1[7:7]);
  C3 I242 (fa3_7min_0[6:6], ct3__0[6:6], termt_2[7:7], termf_1[7:7]);
  C3 I243 (fa3_7min_0[7:7], ct3__0[6:6], termt_2[7:7], termt_1[7:7]);
  NOR3 I244 (simp2361_0[0:0], fa3_7min_0[0:0], fa3_7min_0[3:3], fa3_7min_0[5:5]);
  INV I245 (simp2361_0[1:1], fa3_7min_0[6:6]);
  NAND2 I246 (termf_3[7:7], simp2361_0[0:0], simp2361_0[1:1]);
  NOR3 I247 (simp2371_0[0:0], fa3_7min_0[1:1], fa3_7min_0[2:2], fa3_7min_0[4:4]);
  INV I248 (simp2371_0[1:1], fa3_7min_0[7:7]);
  NAND2 I249 (termt_3[7:7], simp2371_0[0:0], simp2371_0[1:1]);
  AO222 I250 (ct3__0[7:7], termt_1[7:7], termt_2[7:7], termt_1[7:7], ct3__0[6:6], termt_2[7:7], ct3__0[6:6]);
  AO222 I251 (cf3__0[7:7], termf_1[7:7], termf_2[7:7], termf_1[7:7], cf3__0[6:6], termf_2[7:7], cf3__0[6:6]);
  C3 I252 (fa3_8min_0[0:0], cf3__0[7:7], termf_2[8:8], termf_1[8:8]);
  C3 I253 (fa3_8min_0[1:1], cf3__0[7:7], termf_2[8:8], termt_1[8:8]);
  C3 I254 (fa3_8min_0[2:2], cf3__0[7:7], termt_2[8:8], termf_1[8:8]);
  C3 I255 (fa3_8min_0[3:3], cf3__0[7:7], termt_2[8:8], termt_1[8:8]);
  C3 I256 (fa3_8min_0[4:4], ct3__0[7:7], termf_2[8:8], termf_1[8:8]);
  C3 I257 (fa3_8min_0[5:5], ct3__0[7:7], termf_2[8:8], termt_1[8:8]);
  C3 I258 (fa3_8min_0[6:6], ct3__0[7:7], termt_2[8:8], termf_1[8:8]);
  C3 I259 (fa3_8min_0[7:7], ct3__0[7:7], termt_2[8:8], termt_1[8:8]);
  NOR3 I260 (simp2491_0[0:0], fa3_8min_0[0:0], fa3_8min_0[3:3], fa3_8min_0[5:5]);
  INV I261 (simp2491_0[1:1], fa3_8min_0[6:6]);
  NAND2 I262 (termf_3[8:8], simp2491_0[0:0], simp2491_0[1:1]);
  NOR3 I263 (simp2501_0[0:0], fa3_8min_0[1:1], fa3_8min_0[2:2], fa3_8min_0[4:4]);
  INV I264 (simp2501_0[1:1], fa3_8min_0[7:7]);
  NAND2 I265 (termt_3[8:8], simp2501_0[0:0], simp2501_0[1:1]);
  AO222 I266 (ct3__0[8:8], termt_1[8:8], termt_2[8:8], termt_1[8:8], ct3__0[7:7], termt_2[8:8], ct3__0[7:7]);
  AO222 I267 (cf3__0[8:8], termf_1[8:8], termf_2[8:8], termf_1[8:8], cf3__0[7:7], termf_2[8:8], cf3__0[7:7]);
  C3 I268 (fa3_9min_0[0:0], cf3__0[8:8], termf_2[9:9], termf_1[9:9]);
  C3 I269 (fa3_9min_0[1:1], cf3__0[8:8], termf_2[9:9], termt_1[9:9]);
  C3 I270 (fa3_9min_0[2:2], cf3__0[8:8], termt_2[9:9], termf_1[9:9]);
  C3 I271 (fa3_9min_0[3:3], cf3__0[8:8], termt_2[9:9], termt_1[9:9]);
  C3 I272 (fa3_9min_0[4:4], ct3__0[8:8], termf_2[9:9], termf_1[9:9]);
  C3 I273 (fa3_9min_0[5:5], ct3__0[8:8], termf_2[9:9], termt_1[9:9]);
  C3 I274 (fa3_9min_0[6:6], ct3__0[8:8], termt_2[9:9], termf_1[9:9]);
  C3 I275 (fa3_9min_0[7:7], ct3__0[8:8], termt_2[9:9], termt_1[9:9]);
  NOR3 I276 (simp2621_0[0:0], fa3_9min_0[0:0], fa3_9min_0[3:3], fa3_9min_0[5:5]);
  INV I277 (simp2621_0[1:1], fa3_9min_0[6:6]);
  NAND2 I278 (termf_3[9:9], simp2621_0[0:0], simp2621_0[1:1]);
  NOR3 I279 (simp2631_0[0:0], fa3_9min_0[1:1], fa3_9min_0[2:2], fa3_9min_0[4:4]);
  INV I280 (simp2631_0[1:1], fa3_9min_0[7:7]);
  NAND2 I281 (termt_3[9:9], simp2631_0[0:0], simp2631_0[1:1]);
  AO222 I282 (ct3__0[9:9], termt_1[9:9], termt_2[9:9], termt_1[9:9], ct3__0[8:8], termt_2[9:9], ct3__0[8:8]);
  AO222 I283 (cf3__0[9:9], termf_1[9:9], termf_2[9:9], termf_1[9:9], cf3__0[8:8], termf_2[9:9], cf3__0[8:8]);
  C3 I284 (fa3_10min_0[0:0], cf3__0[9:9], termf_2[10:10], termf_1[10:10]);
  C3 I285 (fa3_10min_0[1:1], cf3__0[9:9], termf_2[10:10], termt_1[10:10]);
  C3 I286 (fa3_10min_0[2:2], cf3__0[9:9], termt_2[10:10], termf_1[10:10]);
  C3 I287 (fa3_10min_0[3:3], cf3__0[9:9], termt_2[10:10], termt_1[10:10]);
  C3 I288 (fa3_10min_0[4:4], ct3__0[9:9], termf_2[10:10], termf_1[10:10]);
  C3 I289 (fa3_10min_0[5:5], ct3__0[9:9], termf_2[10:10], termt_1[10:10]);
  C3 I290 (fa3_10min_0[6:6], ct3__0[9:9], termt_2[10:10], termf_1[10:10]);
  C3 I291 (fa3_10min_0[7:7], ct3__0[9:9], termt_2[10:10], termt_1[10:10]);
  NOR3 I292 (simp2751_0[0:0], fa3_10min_0[0:0], fa3_10min_0[3:3], fa3_10min_0[5:5]);
  INV I293 (simp2751_0[1:1], fa3_10min_0[6:6]);
  NAND2 I294 (termf_3[10:10], simp2751_0[0:0], simp2751_0[1:1]);
  NOR3 I295 (simp2761_0[0:0], fa3_10min_0[1:1], fa3_10min_0[2:2], fa3_10min_0[4:4]);
  INV I296 (simp2761_0[1:1], fa3_10min_0[7:7]);
  NAND2 I297 (termt_3[10:10], simp2761_0[0:0], simp2761_0[1:1]);
  AO222 I298 (ct3__0[10:10], termt_1[10:10], termt_2[10:10], termt_1[10:10], ct3__0[9:9], termt_2[10:10], ct3__0[9:9]);
  AO222 I299 (cf3__0[10:10], termf_1[10:10], termf_2[10:10], termf_1[10:10], cf3__0[9:9], termf_2[10:10], cf3__0[9:9]);
  C3 I300 (fa3_11min_0[0:0], cf3__0[10:10], termf_2[11:11], termf_1[11:11]);
  C3 I301 (fa3_11min_0[1:1], cf3__0[10:10], termf_2[11:11], termt_1[11:11]);
  C3 I302 (fa3_11min_0[2:2], cf3__0[10:10], termt_2[11:11], termf_1[11:11]);
  C3 I303 (fa3_11min_0[3:3], cf3__0[10:10], termt_2[11:11], termt_1[11:11]);
  C3 I304 (fa3_11min_0[4:4], ct3__0[10:10], termf_2[11:11], termf_1[11:11]);
  C3 I305 (fa3_11min_0[5:5], ct3__0[10:10], termf_2[11:11], termt_1[11:11]);
  C3 I306 (fa3_11min_0[6:6], ct3__0[10:10], termt_2[11:11], termf_1[11:11]);
  C3 I307 (fa3_11min_0[7:7], ct3__0[10:10], termt_2[11:11], termt_1[11:11]);
  NOR3 I308 (simp2881_0[0:0], fa3_11min_0[0:0], fa3_11min_0[3:3], fa3_11min_0[5:5]);
  INV I309 (simp2881_0[1:1], fa3_11min_0[6:6]);
  NAND2 I310 (termf_3[11:11], simp2881_0[0:0], simp2881_0[1:1]);
  NOR3 I311 (simp2891_0[0:0], fa3_11min_0[1:1], fa3_11min_0[2:2], fa3_11min_0[4:4]);
  INV I312 (simp2891_0[1:1], fa3_11min_0[7:7]);
  NAND2 I313 (termt_3[11:11], simp2891_0[0:0], simp2891_0[1:1]);
  AO222 I314 (ct3__0[11:11], termt_1[11:11], termt_2[11:11], termt_1[11:11], ct3__0[10:10], termt_2[11:11], ct3__0[10:10]);
  AO222 I315 (cf3__0[11:11], termf_1[11:11], termf_2[11:11], termf_1[11:11], cf3__0[10:10], termf_2[11:11], cf3__0[10:10]);
  C3 I316 (fa3_12min_0[0:0], cf3__0[11:11], termf_2[12:12], termf_1[12:12]);
  C3 I317 (fa3_12min_0[1:1], cf3__0[11:11], termf_2[12:12], termt_1[12:12]);
  C3 I318 (fa3_12min_0[2:2], cf3__0[11:11], termt_2[12:12], termf_1[12:12]);
  C3 I319 (fa3_12min_0[3:3], cf3__0[11:11], termt_2[12:12], termt_1[12:12]);
  C3 I320 (fa3_12min_0[4:4], ct3__0[11:11], termf_2[12:12], termf_1[12:12]);
  C3 I321 (fa3_12min_0[5:5], ct3__0[11:11], termf_2[12:12], termt_1[12:12]);
  C3 I322 (fa3_12min_0[6:6], ct3__0[11:11], termt_2[12:12], termf_1[12:12]);
  C3 I323 (fa3_12min_0[7:7], ct3__0[11:11], termt_2[12:12], termt_1[12:12]);
  NOR3 I324 (simp3011_0[0:0], fa3_12min_0[0:0], fa3_12min_0[3:3], fa3_12min_0[5:5]);
  INV I325 (simp3011_0[1:1], fa3_12min_0[6:6]);
  NAND2 I326 (termf_3[12:12], simp3011_0[0:0], simp3011_0[1:1]);
  NOR3 I327 (simp3021_0[0:0], fa3_12min_0[1:1], fa3_12min_0[2:2], fa3_12min_0[4:4]);
  INV I328 (simp3021_0[1:1], fa3_12min_0[7:7]);
  NAND2 I329 (termt_3[12:12], simp3021_0[0:0], simp3021_0[1:1]);
  AO222 I330 (ct3__0[12:12], termt_1[12:12], termt_2[12:12], termt_1[12:12], ct3__0[11:11], termt_2[12:12], ct3__0[11:11]);
  AO222 I331 (cf3__0[12:12], termf_1[12:12], termf_2[12:12], termf_1[12:12], cf3__0[11:11], termf_2[12:12], cf3__0[11:11]);
  C3 I332 (fa3_13min_0[0:0], cf3__0[12:12], termf_2[13:13], termf_1[13:13]);
  C3 I333 (fa3_13min_0[1:1], cf3__0[12:12], termf_2[13:13], termt_1[13:13]);
  C3 I334 (fa3_13min_0[2:2], cf3__0[12:12], termt_2[13:13], termf_1[13:13]);
  C3 I335 (fa3_13min_0[3:3], cf3__0[12:12], termt_2[13:13], termt_1[13:13]);
  C3 I336 (fa3_13min_0[4:4], ct3__0[12:12], termf_2[13:13], termf_1[13:13]);
  C3 I337 (fa3_13min_0[5:5], ct3__0[12:12], termf_2[13:13], termt_1[13:13]);
  C3 I338 (fa3_13min_0[6:6], ct3__0[12:12], termt_2[13:13], termf_1[13:13]);
  C3 I339 (fa3_13min_0[7:7], ct3__0[12:12], termt_2[13:13], termt_1[13:13]);
  NOR3 I340 (simp3141_0[0:0], fa3_13min_0[0:0], fa3_13min_0[3:3], fa3_13min_0[5:5]);
  INV I341 (simp3141_0[1:1], fa3_13min_0[6:6]);
  NAND2 I342 (termf_3[13:13], simp3141_0[0:0], simp3141_0[1:1]);
  NOR3 I343 (simp3151_0[0:0], fa3_13min_0[1:1], fa3_13min_0[2:2], fa3_13min_0[4:4]);
  INV I344 (simp3151_0[1:1], fa3_13min_0[7:7]);
  NAND2 I345 (termt_3[13:13], simp3151_0[0:0], simp3151_0[1:1]);
  AO222 I346 (ct3__0[13:13], termt_1[13:13], termt_2[13:13], termt_1[13:13], ct3__0[12:12], termt_2[13:13], ct3__0[12:12]);
  AO222 I347 (cf3__0[13:13], termf_1[13:13], termf_2[13:13], termf_1[13:13], cf3__0[12:12], termf_2[13:13], cf3__0[12:12]);
  C3 I348 (fa3_14min_0[0:0], cf3__0[13:13], termf_2[14:14], termf_1[14:14]);
  C3 I349 (fa3_14min_0[1:1], cf3__0[13:13], termf_2[14:14], termt_1[14:14]);
  C3 I350 (fa3_14min_0[2:2], cf3__0[13:13], termt_2[14:14], termf_1[14:14]);
  C3 I351 (fa3_14min_0[3:3], cf3__0[13:13], termt_2[14:14], termt_1[14:14]);
  C3 I352 (fa3_14min_0[4:4], ct3__0[13:13], termf_2[14:14], termf_1[14:14]);
  C3 I353 (fa3_14min_0[5:5], ct3__0[13:13], termf_2[14:14], termt_1[14:14]);
  C3 I354 (fa3_14min_0[6:6], ct3__0[13:13], termt_2[14:14], termf_1[14:14]);
  C3 I355 (fa3_14min_0[7:7], ct3__0[13:13], termt_2[14:14], termt_1[14:14]);
  NOR3 I356 (simp3271_0[0:0], fa3_14min_0[0:0], fa3_14min_0[3:3], fa3_14min_0[5:5]);
  INV I357 (simp3271_0[1:1], fa3_14min_0[6:6]);
  NAND2 I358 (termf_3[14:14], simp3271_0[0:0], simp3271_0[1:1]);
  NOR3 I359 (simp3281_0[0:0], fa3_14min_0[1:1], fa3_14min_0[2:2], fa3_14min_0[4:4]);
  INV I360 (simp3281_0[1:1], fa3_14min_0[7:7]);
  NAND2 I361 (termt_3[14:14], simp3281_0[0:0], simp3281_0[1:1]);
  AO222 I362 (ct3__0[14:14], termt_1[14:14], termt_2[14:14], termt_1[14:14], ct3__0[13:13], termt_2[14:14], ct3__0[13:13]);
  AO222 I363 (cf3__0[14:14], termf_1[14:14], termf_2[14:14], termf_1[14:14], cf3__0[13:13], termf_2[14:14], cf3__0[13:13]);
  C3 I364 (fa3_15min_0[0:0], cf3__0[14:14], termf_2[15:15], termf_1[15:15]);
  C3 I365 (fa3_15min_0[1:1], cf3__0[14:14], termf_2[15:15], termt_1[15:15]);
  C3 I366 (fa3_15min_0[2:2], cf3__0[14:14], termt_2[15:15], termf_1[15:15]);
  C3 I367 (fa3_15min_0[3:3], cf3__0[14:14], termt_2[15:15], termt_1[15:15]);
  C3 I368 (fa3_15min_0[4:4], ct3__0[14:14], termf_2[15:15], termf_1[15:15]);
  C3 I369 (fa3_15min_0[5:5], ct3__0[14:14], termf_2[15:15], termt_1[15:15]);
  C3 I370 (fa3_15min_0[6:6], ct3__0[14:14], termt_2[15:15], termf_1[15:15]);
  C3 I371 (fa3_15min_0[7:7], ct3__0[14:14], termt_2[15:15], termt_1[15:15]);
  NOR3 I372 (simp3401_0[0:0], fa3_15min_0[0:0], fa3_15min_0[3:3], fa3_15min_0[5:5]);
  INV I373 (simp3401_0[1:1], fa3_15min_0[6:6]);
  NAND2 I374 (termf_3[15:15], simp3401_0[0:0], simp3401_0[1:1]);
  NOR3 I375 (simp3411_0[0:0], fa3_15min_0[1:1], fa3_15min_0[2:2], fa3_15min_0[4:4]);
  INV I376 (simp3411_0[1:1], fa3_15min_0[7:7]);
  NAND2 I377 (termt_3[15:15], simp3411_0[0:0], simp3411_0[1:1]);
  AO222 I378 (ct3__0[15:15], termt_1[15:15], termt_2[15:15], termt_1[15:15], ct3__0[14:14], termt_2[15:15], ct3__0[14:14]);
  AO222 I379 (cf3__0[15:15], termf_1[15:15], termf_2[15:15], termf_1[15:15], cf3__0[14:14], termf_2[15:15], cf3__0[14:14]);
  C3 I380 (fa3_16min_0[0:0], cf3__0[15:15], termf_2[16:16], termf_1[16:16]);
  C3 I381 (fa3_16min_0[1:1], cf3__0[15:15], termf_2[16:16], termt_1[16:16]);
  C3 I382 (fa3_16min_0[2:2], cf3__0[15:15], termt_2[16:16], termf_1[16:16]);
  C3 I383 (fa3_16min_0[3:3], cf3__0[15:15], termt_2[16:16], termt_1[16:16]);
  C3 I384 (fa3_16min_0[4:4], ct3__0[15:15], termf_2[16:16], termf_1[16:16]);
  C3 I385 (fa3_16min_0[5:5], ct3__0[15:15], termf_2[16:16], termt_1[16:16]);
  C3 I386 (fa3_16min_0[6:6], ct3__0[15:15], termt_2[16:16], termf_1[16:16]);
  C3 I387 (fa3_16min_0[7:7], ct3__0[15:15], termt_2[16:16], termt_1[16:16]);
  NOR3 I388 (simp3531_0[0:0], fa3_16min_0[0:0], fa3_16min_0[3:3], fa3_16min_0[5:5]);
  INV I389 (simp3531_0[1:1], fa3_16min_0[6:6]);
  NAND2 I390 (termf_3[16:16], simp3531_0[0:0], simp3531_0[1:1]);
  NOR3 I391 (simp3541_0[0:0], fa3_16min_0[1:1], fa3_16min_0[2:2], fa3_16min_0[4:4]);
  INV I392 (simp3541_0[1:1], fa3_16min_0[7:7]);
  NAND2 I393 (termt_3[16:16], simp3541_0[0:0], simp3541_0[1:1]);
  AO222 I394 (ct3__0[16:16], termt_1[16:16], termt_2[16:16], termt_1[16:16], ct3__0[15:15], termt_2[16:16], ct3__0[15:15]);
  AO222 I395 (cf3__0[16:16], termf_1[16:16], termf_2[16:16], termf_1[16:16], cf3__0[15:15], termf_2[16:16], cf3__0[15:15]);
  C3 I396 (fa3_17min_0[0:0], cf3__0[16:16], termf_2[17:17], termf_1[17:17]);
  C3 I397 (fa3_17min_0[1:1], cf3__0[16:16], termf_2[17:17], termt_1[17:17]);
  C3 I398 (fa3_17min_0[2:2], cf3__0[16:16], termt_2[17:17], termf_1[17:17]);
  C3 I399 (fa3_17min_0[3:3], cf3__0[16:16], termt_2[17:17], termt_1[17:17]);
  C3 I400 (fa3_17min_0[4:4], ct3__0[16:16], termf_2[17:17], termf_1[17:17]);
  C3 I401 (fa3_17min_0[5:5], ct3__0[16:16], termf_2[17:17], termt_1[17:17]);
  C3 I402 (fa3_17min_0[6:6], ct3__0[16:16], termt_2[17:17], termf_1[17:17]);
  C3 I403 (fa3_17min_0[7:7], ct3__0[16:16], termt_2[17:17], termt_1[17:17]);
  NOR3 I404 (simp3661_0[0:0], fa3_17min_0[0:0], fa3_17min_0[3:3], fa3_17min_0[5:5]);
  INV I405 (simp3661_0[1:1], fa3_17min_0[6:6]);
  NAND2 I406 (termf_3[17:17], simp3661_0[0:0], simp3661_0[1:1]);
  NOR3 I407 (simp3671_0[0:0], fa3_17min_0[1:1], fa3_17min_0[2:2], fa3_17min_0[4:4]);
  INV I408 (simp3671_0[1:1], fa3_17min_0[7:7]);
  NAND2 I409 (termt_3[17:17], simp3671_0[0:0], simp3671_0[1:1]);
  AO222 I410 (ct3__0[17:17], termt_1[17:17], termt_2[17:17], termt_1[17:17], ct3__0[16:16], termt_2[17:17], ct3__0[16:16]);
  AO222 I411 (cf3__0[17:17], termf_1[17:17], termf_2[17:17], termf_1[17:17], cf3__0[16:16], termf_2[17:17], cf3__0[16:16]);
  C3 I412 (fa3_18min_0[0:0], cf3__0[17:17], termf_2[18:18], termf_1[18:18]);
  C3 I413 (fa3_18min_0[1:1], cf3__0[17:17], termf_2[18:18], termt_1[18:18]);
  C3 I414 (fa3_18min_0[2:2], cf3__0[17:17], termt_2[18:18], termf_1[18:18]);
  C3 I415 (fa3_18min_0[3:3], cf3__0[17:17], termt_2[18:18], termt_1[18:18]);
  C3 I416 (fa3_18min_0[4:4], ct3__0[17:17], termf_2[18:18], termf_1[18:18]);
  C3 I417 (fa3_18min_0[5:5], ct3__0[17:17], termf_2[18:18], termt_1[18:18]);
  C3 I418 (fa3_18min_0[6:6], ct3__0[17:17], termt_2[18:18], termf_1[18:18]);
  C3 I419 (fa3_18min_0[7:7], ct3__0[17:17], termt_2[18:18], termt_1[18:18]);
  NOR3 I420 (simp3791_0[0:0], fa3_18min_0[0:0], fa3_18min_0[3:3], fa3_18min_0[5:5]);
  INV I421 (simp3791_0[1:1], fa3_18min_0[6:6]);
  NAND2 I422 (termf_3[18:18], simp3791_0[0:0], simp3791_0[1:1]);
  NOR3 I423 (simp3801_0[0:0], fa3_18min_0[1:1], fa3_18min_0[2:2], fa3_18min_0[4:4]);
  INV I424 (simp3801_0[1:1], fa3_18min_0[7:7]);
  NAND2 I425 (termt_3[18:18], simp3801_0[0:0], simp3801_0[1:1]);
  AO222 I426 (ct3__0[18:18], termt_1[18:18], termt_2[18:18], termt_1[18:18], ct3__0[17:17], termt_2[18:18], ct3__0[17:17]);
  AO222 I427 (cf3__0[18:18], termf_1[18:18], termf_2[18:18], termf_1[18:18], cf3__0[17:17], termf_2[18:18], cf3__0[17:17]);
  C3 I428 (fa3_19min_0[0:0], cf3__0[18:18], termf_2[19:19], termf_1[19:19]);
  C3 I429 (fa3_19min_0[1:1], cf3__0[18:18], termf_2[19:19], termt_1[19:19]);
  C3 I430 (fa3_19min_0[2:2], cf3__0[18:18], termt_2[19:19], termf_1[19:19]);
  C3 I431 (fa3_19min_0[3:3], cf3__0[18:18], termt_2[19:19], termt_1[19:19]);
  C3 I432 (fa3_19min_0[4:4], ct3__0[18:18], termf_2[19:19], termf_1[19:19]);
  C3 I433 (fa3_19min_0[5:5], ct3__0[18:18], termf_2[19:19], termt_1[19:19]);
  C3 I434 (fa3_19min_0[6:6], ct3__0[18:18], termt_2[19:19], termf_1[19:19]);
  C3 I435 (fa3_19min_0[7:7], ct3__0[18:18], termt_2[19:19], termt_1[19:19]);
  NOR3 I436 (simp3921_0[0:0], fa3_19min_0[0:0], fa3_19min_0[3:3], fa3_19min_0[5:5]);
  INV I437 (simp3921_0[1:1], fa3_19min_0[6:6]);
  NAND2 I438 (termf_3[19:19], simp3921_0[0:0], simp3921_0[1:1]);
  NOR3 I439 (simp3931_0[0:0], fa3_19min_0[1:1], fa3_19min_0[2:2], fa3_19min_0[4:4]);
  INV I440 (simp3931_0[1:1], fa3_19min_0[7:7]);
  NAND2 I441 (termt_3[19:19], simp3931_0[0:0], simp3931_0[1:1]);
  AO222 I442 (ct3__0[19:19], termt_1[19:19], termt_2[19:19], termt_1[19:19], ct3__0[18:18], termt_2[19:19], ct3__0[18:18]);
  AO222 I443 (cf3__0[19:19], termf_1[19:19], termf_2[19:19], termf_1[19:19], cf3__0[18:18], termf_2[19:19], cf3__0[18:18]);
  C3 I444 (fa3_20min_0[0:0], cf3__0[19:19], termf_2[20:20], termf_1[20:20]);
  C3 I445 (fa3_20min_0[1:1], cf3__0[19:19], termf_2[20:20], termt_1[20:20]);
  C3 I446 (fa3_20min_0[2:2], cf3__0[19:19], termt_2[20:20], termf_1[20:20]);
  C3 I447 (fa3_20min_0[3:3], cf3__0[19:19], termt_2[20:20], termt_1[20:20]);
  C3 I448 (fa3_20min_0[4:4], ct3__0[19:19], termf_2[20:20], termf_1[20:20]);
  C3 I449 (fa3_20min_0[5:5], ct3__0[19:19], termf_2[20:20], termt_1[20:20]);
  C3 I450 (fa3_20min_0[6:6], ct3__0[19:19], termt_2[20:20], termf_1[20:20]);
  C3 I451 (fa3_20min_0[7:7], ct3__0[19:19], termt_2[20:20], termt_1[20:20]);
  NOR3 I452 (simp4051_0[0:0], fa3_20min_0[0:0], fa3_20min_0[3:3], fa3_20min_0[5:5]);
  INV I453 (simp4051_0[1:1], fa3_20min_0[6:6]);
  NAND2 I454 (termf_3[20:20], simp4051_0[0:0], simp4051_0[1:1]);
  NOR3 I455 (simp4061_0[0:0], fa3_20min_0[1:1], fa3_20min_0[2:2], fa3_20min_0[4:4]);
  INV I456 (simp4061_0[1:1], fa3_20min_0[7:7]);
  NAND2 I457 (termt_3[20:20], simp4061_0[0:0], simp4061_0[1:1]);
  AO222 I458 (ct3__0[20:20], termt_1[20:20], termt_2[20:20], termt_1[20:20], ct3__0[19:19], termt_2[20:20], ct3__0[19:19]);
  AO222 I459 (cf3__0[20:20], termf_1[20:20], termf_2[20:20], termf_1[20:20], cf3__0[19:19], termf_2[20:20], cf3__0[19:19]);
  C3 I460 (fa3_21min_0[0:0], cf3__0[20:20], termf_2[21:21], termf_1[21:21]);
  C3 I461 (fa3_21min_0[1:1], cf3__0[20:20], termf_2[21:21], termt_1[21:21]);
  C3 I462 (fa3_21min_0[2:2], cf3__0[20:20], termt_2[21:21], termf_1[21:21]);
  C3 I463 (fa3_21min_0[3:3], cf3__0[20:20], termt_2[21:21], termt_1[21:21]);
  C3 I464 (fa3_21min_0[4:4], ct3__0[20:20], termf_2[21:21], termf_1[21:21]);
  C3 I465 (fa3_21min_0[5:5], ct3__0[20:20], termf_2[21:21], termt_1[21:21]);
  C3 I466 (fa3_21min_0[6:6], ct3__0[20:20], termt_2[21:21], termf_1[21:21]);
  C3 I467 (fa3_21min_0[7:7], ct3__0[20:20], termt_2[21:21], termt_1[21:21]);
  NOR3 I468 (simp4181_0[0:0], fa3_21min_0[0:0], fa3_21min_0[3:3], fa3_21min_0[5:5]);
  INV I469 (simp4181_0[1:1], fa3_21min_0[6:6]);
  NAND2 I470 (termf_3[21:21], simp4181_0[0:0], simp4181_0[1:1]);
  NOR3 I471 (simp4191_0[0:0], fa3_21min_0[1:1], fa3_21min_0[2:2], fa3_21min_0[4:4]);
  INV I472 (simp4191_0[1:1], fa3_21min_0[7:7]);
  NAND2 I473 (termt_3[21:21], simp4191_0[0:0], simp4191_0[1:1]);
  AO222 I474 (ct3__0[21:21], termt_1[21:21], termt_2[21:21], termt_1[21:21], ct3__0[20:20], termt_2[21:21], ct3__0[20:20]);
  AO222 I475 (cf3__0[21:21], termf_1[21:21], termf_2[21:21], termf_1[21:21], cf3__0[20:20], termf_2[21:21], cf3__0[20:20]);
  C3 I476 (fa3_22min_0[0:0], cf3__0[21:21], termf_2[22:22], termf_1[22:22]);
  C3 I477 (fa3_22min_0[1:1], cf3__0[21:21], termf_2[22:22], termt_1[22:22]);
  C3 I478 (fa3_22min_0[2:2], cf3__0[21:21], termt_2[22:22], termf_1[22:22]);
  C3 I479 (fa3_22min_0[3:3], cf3__0[21:21], termt_2[22:22], termt_1[22:22]);
  C3 I480 (fa3_22min_0[4:4], ct3__0[21:21], termf_2[22:22], termf_1[22:22]);
  C3 I481 (fa3_22min_0[5:5], ct3__0[21:21], termf_2[22:22], termt_1[22:22]);
  C3 I482 (fa3_22min_0[6:6], ct3__0[21:21], termt_2[22:22], termf_1[22:22]);
  C3 I483 (fa3_22min_0[7:7], ct3__0[21:21], termt_2[22:22], termt_1[22:22]);
  NOR3 I484 (simp4311_0[0:0], fa3_22min_0[0:0], fa3_22min_0[3:3], fa3_22min_0[5:5]);
  INV I485 (simp4311_0[1:1], fa3_22min_0[6:6]);
  NAND2 I486 (termf_3[22:22], simp4311_0[0:0], simp4311_0[1:1]);
  NOR3 I487 (simp4321_0[0:0], fa3_22min_0[1:1], fa3_22min_0[2:2], fa3_22min_0[4:4]);
  INV I488 (simp4321_0[1:1], fa3_22min_0[7:7]);
  NAND2 I489 (termt_3[22:22], simp4321_0[0:0], simp4321_0[1:1]);
  AO222 I490 (ct3__0[22:22], termt_1[22:22], termt_2[22:22], termt_1[22:22], ct3__0[21:21], termt_2[22:22], ct3__0[21:21]);
  AO222 I491 (cf3__0[22:22], termf_1[22:22], termf_2[22:22], termf_1[22:22], cf3__0[21:21], termf_2[22:22], cf3__0[21:21]);
  C3 I492 (fa3_23min_0[0:0], cf3__0[22:22], termf_2[23:23], termf_1[23:23]);
  C3 I493 (fa3_23min_0[1:1], cf3__0[22:22], termf_2[23:23], termt_1[23:23]);
  C3 I494 (fa3_23min_0[2:2], cf3__0[22:22], termt_2[23:23], termf_1[23:23]);
  C3 I495 (fa3_23min_0[3:3], cf3__0[22:22], termt_2[23:23], termt_1[23:23]);
  C3 I496 (fa3_23min_0[4:4], ct3__0[22:22], termf_2[23:23], termf_1[23:23]);
  C3 I497 (fa3_23min_0[5:5], ct3__0[22:22], termf_2[23:23], termt_1[23:23]);
  C3 I498 (fa3_23min_0[6:6], ct3__0[22:22], termt_2[23:23], termf_1[23:23]);
  C3 I499 (fa3_23min_0[7:7], ct3__0[22:22], termt_2[23:23], termt_1[23:23]);
  NOR3 I500 (simp4441_0[0:0], fa3_23min_0[0:0], fa3_23min_0[3:3], fa3_23min_0[5:5]);
  INV I501 (simp4441_0[1:1], fa3_23min_0[6:6]);
  NAND2 I502 (termf_3[23:23], simp4441_0[0:0], simp4441_0[1:1]);
  NOR3 I503 (simp4451_0[0:0], fa3_23min_0[1:1], fa3_23min_0[2:2], fa3_23min_0[4:4]);
  INV I504 (simp4451_0[1:1], fa3_23min_0[7:7]);
  NAND2 I505 (termt_3[23:23], simp4451_0[0:0], simp4451_0[1:1]);
  AO222 I506 (ct3__0[23:23], termt_1[23:23], termt_2[23:23], termt_1[23:23], ct3__0[22:22], termt_2[23:23], ct3__0[22:22]);
  AO222 I507 (cf3__0[23:23], termf_1[23:23], termf_2[23:23], termf_1[23:23], cf3__0[22:22], termf_2[23:23], cf3__0[22:22]);
  C3 I508 (fa3_24min_0[0:0], cf3__0[23:23], termf_2[24:24], termf_1[24:24]);
  C3 I509 (fa3_24min_0[1:1], cf3__0[23:23], termf_2[24:24], termt_1[24:24]);
  C3 I510 (fa3_24min_0[2:2], cf3__0[23:23], termt_2[24:24], termf_1[24:24]);
  C3 I511 (fa3_24min_0[3:3], cf3__0[23:23], termt_2[24:24], termt_1[24:24]);
  C3 I512 (fa3_24min_0[4:4], ct3__0[23:23], termf_2[24:24], termf_1[24:24]);
  C3 I513 (fa3_24min_0[5:5], ct3__0[23:23], termf_2[24:24], termt_1[24:24]);
  C3 I514 (fa3_24min_0[6:6], ct3__0[23:23], termt_2[24:24], termf_1[24:24]);
  C3 I515 (fa3_24min_0[7:7], ct3__0[23:23], termt_2[24:24], termt_1[24:24]);
  NOR3 I516 (simp4571_0[0:0], fa3_24min_0[0:0], fa3_24min_0[3:3], fa3_24min_0[5:5]);
  INV I517 (simp4571_0[1:1], fa3_24min_0[6:6]);
  NAND2 I518 (termf_3[24:24], simp4571_0[0:0], simp4571_0[1:1]);
  NOR3 I519 (simp4581_0[0:0], fa3_24min_0[1:1], fa3_24min_0[2:2], fa3_24min_0[4:4]);
  INV I520 (simp4581_0[1:1], fa3_24min_0[7:7]);
  NAND2 I521 (termt_3[24:24], simp4581_0[0:0], simp4581_0[1:1]);
  AO222 I522 (ct3__0[24:24], termt_1[24:24], termt_2[24:24], termt_1[24:24], ct3__0[23:23], termt_2[24:24], ct3__0[23:23]);
  AO222 I523 (cf3__0[24:24], termf_1[24:24], termf_2[24:24], termf_1[24:24], cf3__0[23:23], termf_2[24:24], cf3__0[23:23]);
  C3 I524 (fa3_25min_0[0:0], cf3__0[24:24], termf_2[25:25], termf_1[25:25]);
  C3 I525 (fa3_25min_0[1:1], cf3__0[24:24], termf_2[25:25], termt_1[25:25]);
  C3 I526 (fa3_25min_0[2:2], cf3__0[24:24], termt_2[25:25], termf_1[25:25]);
  C3 I527 (fa3_25min_0[3:3], cf3__0[24:24], termt_2[25:25], termt_1[25:25]);
  C3 I528 (fa3_25min_0[4:4], ct3__0[24:24], termf_2[25:25], termf_1[25:25]);
  C3 I529 (fa3_25min_0[5:5], ct3__0[24:24], termf_2[25:25], termt_1[25:25]);
  C3 I530 (fa3_25min_0[6:6], ct3__0[24:24], termt_2[25:25], termf_1[25:25]);
  C3 I531 (fa3_25min_0[7:7], ct3__0[24:24], termt_2[25:25], termt_1[25:25]);
  NOR3 I532 (simp4701_0[0:0], fa3_25min_0[0:0], fa3_25min_0[3:3], fa3_25min_0[5:5]);
  INV I533 (simp4701_0[1:1], fa3_25min_0[6:6]);
  NAND2 I534 (termf_3[25:25], simp4701_0[0:0], simp4701_0[1:1]);
  NOR3 I535 (simp4711_0[0:0], fa3_25min_0[1:1], fa3_25min_0[2:2], fa3_25min_0[4:4]);
  INV I536 (simp4711_0[1:1], fa3_25min_0[7:7]);
  NAND2 I537 (termt_3[25:25], simp4711_0[0:0], simp4711_0[1:1]);
  AO222 I538 (ct3__0[25:25], termt_1[25:25], termt_2[25:25], termt_1[25:25], ct3__0[24:24], termt_2[25:25], ct3__0[24:24]);
  AO222 I539 (cf3__0[25:25], termf_1[25:25], termf_2[25:25], termf_1[25:25], cf3__0[24:24], termf_2[25:25], cf3__0[24:24]);
  C3 I540 (fa3_26min_0[0:0], cf3__0[25:25], termf_2[26:26], termf_1[26:26]);
  C3 I541 (fa3_26min_0[1:1], cf3__0[25:25], termf_2[26:26], termt_1[26:26]);
  C3 I542 (fa3_26min_0[2:2], cf3__0[25:25], termt_2[26:26], termf_1[26:26]);
  C3 I543 (fa3_26min_0[3:3], cf3__0[25:25], termt_2[26:26], termt_1[26:26]);
  C3 I544 (fa3_26min_0[4:4], ct3__0[25:25], termf_2[26:26], termf_1[26:26]);
  C3 I545 (fa3_26min_0[5:5], ct3__0[25:25], termf_2[26:26], termt_1[26:26]);
  C3 I546 (fa3_26min_0[6:6], ct3__0[25:25], termt_2[26:26], termf_1[26:26]);
  C3 I547 (fa3_26min_0[7:7], ct3__0[25:25], termt_2[26:26], termt_1[26:26]);
  NOR3 I548 (simp4831_0[0:0], fa3_26min_0[0:0], fa3_26min_0[3:3], fa3_26min_0[5:5]);
  INV I549 (simp4831_0[1:1], fa3_26min_0[6:6]);
  NAND2 I550 (termf_3[26:26], simp4831_0[0:0], simp4831_0[1:1]);
  NOR3 I551 (simp4841_0[0:0], fa3_26min_0[1:1], fa3_26min_0[2:2], fa3_26min_0[4:4]);
  INV I552 (simp4841_0[1:1], fa3_26min_0[7:7]);
  NAND2 I553 (termt_3[26:26], simp4841_0[0:0], simp4841_0[1:1]);
  AO222 I554 (ct3__0[26:26], termt_1[26:26], termt_2[26:26], termt_1[26:26], ct3__0[25:25], termt_2[26:26], ct3__0[25:25]);
  AO222 I555 (cf3__0[26:26], termf_1[26:26], termf_2[26:26], termf_1[26:26], cf3__0[25:25], termf_2[26:26], cf3__0[25:25]);
  C3 I556 (fa3_27min_0[0:0], cf3__0[26:26], termf_2[27:27], termf_1[27:27]);
  C3 I557 (fa3_27min_0[1:1], cf3__0[26:26], termf_2[27:27], termt_1[27:27]);
  C3 I558 (fa3_27min_0[2:2], cf3__0[26:26], termt_2[27:27], termf_1[27:27]);
  C3 I559 (fa3_27min_0[3:3], cf3__0[26:26], termt_2[27:27], termt_1[27:27]);
  C3 I560 (fa3_27min_0[4:4], ct3__0[26:26], termf_2[27:27], termf_1[27:27]);
  C3 I561 (fa3_27min_0[5:5], ct3__0[26:26], termf_2[27:27], termt_1[27:27]);
  C3 I562 (fa3_27min_0[6:6], ct3__0[26:26], termt_2[27:27], termf_1[27:27]);
  C3 I563 (fa3_27min_0[7:7], ct3__0[26:26], termt_2[27:27], termt_1[27:27]);
  NOR3 I564 (simp4961_0[0:0], fa3_27min_0[0:0], fa3_27min_0[3:3], fa3_27min_0[5:5]);
  INV I565 (simp4961_0[1:1], fa3_27min_0[6:6]);
  NAND2 I566 (termf_3[27:27], simp4961_0[0:0], simp4961_0[1:1]);
  NOR3 I567 (simp4971_0[0:0], fa3_27min_0[1:1], fa3_27min_0[2:2], fa3_27min_0[4:4]);
  INV I568 (simp4971_0[1:1], fa3_27min_0[7:7]);
  NAND2 I569 (termt_3[27:27], simp4971_0[0:0], simp4971_0[1:1]);
  AO222 I570 (ct3__0[27:27], termt_1[27:27], termt_2[27:27], termt_1[27:27], ct3__0[26:26], termt_2[27:27], ct3__0[26:26]);
  AO222 I571 (cf3__0[27:27], termf_1[27:27], termf_2[27:27], termf_1[27:27], cf3__0[26:26], termf_2[27:27], cf3__0[26:26]);
  C3 I572 (fa3_28min_0[0:0], cf3__0[27:27], termf_2[28:28], termf_1[28:28]);
  C3 I573 (fa3_28min_0[1:1], cf3__0[27:27], termf_2[28:28], termt_1[28:28]);
  C3 I574 (fa3_28min_0[2:2], cf3__0[27:27], termt_2[28:28], termf_1[28:28]);
  C3 I575 (fa3_28min_0[3:3], cf3__0[27:27], termt_2[28:28], termt_1[28:28]);
  C3 I576 (fa3_28min_0[4:4], ct3__0[27:27], termf_2[28:28], termf_1[28:28]);
  C3 I577 (fa3_28min_0[5:5], ct3__0[27:27], termf_2[28:28], termt_1[28:28]);
  C3 I578 (fa3_28min_0[6:6], ct3__0[27:27], termt_2[28:28], termf_1[28:28]);
  C3 I579 (fa3_28min_0[7:7], ct3__0[27:27], termt_2[28:28], termt_1[28:28]);
  NOR3 I580 (simp5091_0[0:0], fa3_28min_0[0:0], fa3_28min_0[3:3], fa3_28min_0[5:5]);
  INV I581 (simp5091_0[1:1], fa3_28min_0[6:6]);
  NAND2 I582 (termf_3[28:28], simp5091_0[0:0], simp5091_0[1:1]);
  NOR3 I583 (simp5101_0[0:0], fa3_28min_0[1:1], fa3_28min_0[2:2], fa3_28min_0[4:4]);
  INV I584 (simp5101_0[1:1], fa3_28min_0[7:7]);
  NAND2 I585 (termt_3[28:28], simp5101_0[0:0], simp5101_0[1:1]);
  AO222 I586 (ct3__0[28:28], termt_1[28:28], termt_2[28:28], termt_1[28:28], ct3__0[27:27], termt_2[28:28], ct3__0[27:27]);
  AO222 I587 (cf3__0[28:28], termf_1[28:28], termf_2[28:28], termf_1[28:28], cf3__0[27:27], termf_2[28:28], cf3__0[27:27]);
  C3 I588 (fa3_29min_0[0:0], cf3__0[28:28], termf_2[29:29], termf_1[29:29]);
  C3 I589 (fa3_29min_0[1:1], cf3__0[28:28], termf_2[29:29], termt_1[29:29]);
  C3 I590 (fa3_29min_0[2:2], cf3__0[28:28], termt_2[29:29], termf_1[29:29]);
  C3 I591 (fa3_29min_0[3:3], cf3__0[28:28], termt_2[29:29], termt_1[29:29]);
  C3 I592 (fa3_29min_0[4:4], ct3__0[28:28], termf_2[29:29], termf_1[29:29]);
  C3 I593 (fa3_29min_0[5:5], ct3__0[28:28], termf_2[29:29], termt_1[29:29]);
  C3 I594 (fa3_29min_0[6:6], ct3__0[28:28], termt_2[29:29], termf_1[29:29]);
  C3 I595 (fa3_29min_0[7:7], ct3__0[28:28], termt_2[29:29], termt_1[29:29]);
  NOR3 I596 (simp5221_0[0:0], fa3_29min_0[0:0], fa3_29min_0[3:3], fa3_29min_0[5:5]);
  INV I597 (simp5221_0[1:1], fa3_29min_0[6:6]);
  NAND2 I598 (termf_3[29:29], simp5221_0[0:0], simp5221_0[1:1]);
  NOR3 I599 (simp5231_0[0:0], fa3_29min_0[1:1], fa3_29min_0[2:2], fa3_29min_0[4:4]);
  INV I600 (simp5231_0[1:1], fa3_29min_0[7:7]);
  NAND2 I601 (termt_3[29:29], simp5231_0[0:0], simp5231_0[1:1]);
  AO222 I602 (ct3__0[29:29], termt_1[29:29], termt_2[29:29], termt_1[29:29], ct3__0[28:28], termt_2[29:29], ct3__0[28:28]);
  AO222 I603 (cf3__0[29:29], termf_1[29:29], termf_2[29:29], termf_1[29:29], cf3__0[28:28], termf_2[29:29], cf3__0[28:28]);
  C3 I604 (fa3_30min_0[0:0], cf3__0[29:29], termf_2[30:30], termf_1[30:30]);
  C3 I605 (fa3_30min_0[1:1], cf3__0[29:29], termf_2[30:30], termt_1[30:30]);
  C3 I606 (fa3_30min_0[2:2], cf3__0[29:29], termt_2[30:30], termf_1[30:30]);
  C3 I607 (fa3_30min_0[3:3], cf3__0[29:29], termt_2[30:30], termt_1[30:30]);
  C3 I608 (fa3_30min_0[4:4], ct3__0[29:29], termf_2[30:30], termf_1[30:30]);
  C3 I609 (fa3_30min_0[5:5], ct3__0[29:29], termf_2[30:30], termt_1[30:30]);
  C3 I610 (fa3_30min_0[6:6], ct3__0[29:29], termt_2[30:30], termf_1[30:30]);
  C3 I611 (fa3_30min_0[7:7], ct3__0[29:29], termt_2[30:30], termt_1[30:30]);
  NOR3 I612 (simp5351_0[0:0], fa3_30min_0[0:0], fa3_30min_0[3:3], fa3_30min_0[5:5]);
  INV I613 (simp5351_0[1:1], fa3_30min_0[6:6]);
  NAND2 I614 (termf_3[30:30], simp5351_0[0:0], simp5351_0[1:1]);
  NOR3 I615 (simp5361_0[0:0], fa3_30min_0[1:1], fa3_30min_0[2:2], fa3_30min_0[4:4]);
  INV I616 (simp5361_0[1:1], fa3_30min_0[7:7]);
  NAND2 I617 (termt_3[30:30], simp5361_0[0:0], simp5361_0[1:1]);
  AO222 I618 (ct3__0[30:30], termt_1[30:30], termt_2[30:30], termt_1[30:30], ct3__0[29:29], termt_2[30:30], ct3__0[29:29]);
  AO222 I619 (cf3__0[30:30], termf_1[30:30], termf_2[30:30], termf_1[30:30], cf3__0[29:29], termf_2[30:30], cf3__0[29:29]);
  C3 I620 (fa3_31min_0[0:0], cf3__0[30:30], termf_2[31:31], termf_1[31:31]);
  C3 I621 (fa3_31min_0[1:1], cf3__0[30:30], termf_2[31:31], termt_1[31:31]);
  C3 I622 (fa3_31min_0[2:2], cf3__0[30:30], termt_2[31:31], termf_1[31:31]);
  C3 I623 (fa3_31min_0[3:3], cf3__0[30:30], termt_2[31:31], termt_1[31:31]);
  C3 I624 (fa3_31min_0[4:4], ct3__0[30:30], termf_2[31:31], termf_1[31:31]);
  C3 I625 (fa3_31min_0[5:5], ct3__0[30:30], termf_2[31:31], termt_1[31:31]);
  C3 I626 (fa3_31min_0[6:6], ct3__0[30:30], termt_2[31:31], termf_1[31:31]);
  C3 I627 (fa3_31min_0[7:7], ct3__0[30:30], termt_2[31:31], termt_1[31:31]);
  NOR3 I628 (simp5481_0[0:0], fa3_31min_0[0:0], fa3_31min_0[3:3], fa3_31min_0[5:5]);
  INV I629 (simp5481_0[1:1], fa3_31min_0[6:6]);
  NAND2 I630 (termf_3[31:31], simp5481_0[0:0], simp5481_0[1:1]);
  NOR3 I631 (simp5491_0[0:0], fa3_31min_0[1:1], fa3_31min_0[2:2], fa3_31min_0[4:4]);
  INV I632 (simp5491_0[1:1], fa3_31min_0[7:7]);
  NAND2 I633 (termt_3[31:31], simp5491_0[0:0], simp5491_0[1:1]);
  AO222 I634 (ct3__0[31:31], termt_1[31:31], termt_2[31:31], termt_1[31:31], ct3__0[30:30], termt_2[31:31], ct3__0[30:30]);
  AO222 I635 (cf3__0[31:31], termf_1[31:31], termf_2[31:31], termf_1[31:31], cf3__0[30:30], termf_2[31:31], cf3__0[30:30]);
  C3 I636 (fa3_32min_0[0:0], cf3__0[31:31], termf_2[32:32], termf_1[32:32]);
  C3 I637 (fa3_32min_0[1:1], cf3__0[31:31], termf_2[32:32], termt_1[32:32]);
  C3 I638 (fa3_32min_0[2:2], cf3__0[31:31], termt_2[32:32], termf_1[32:32]);
  C3 I639 (fa3_32min_0[3:3], cf3__0[31:31], termt_2[32:32], termt_1[32:32]);
  C3 I640 (fa3_32min_0[4:4], ct3__0[31:31], termf_2[32:32], termf_1[32:32]);
  C3 I641 (fa3_32min_0[5:5], ct3__0[31:31], termf_2[32:32], termt_1[32:32]);
  C3 I642 (fa3_32min_0[6:6], ct3__0[31:31], termt_2[32:32], termf_1[32:32]);
  C3 I643 (fa3_32min_0[7:7], ct3__0[31:31], termt_2[32:32], termt_1[32:32]);
  NOR3 I644 (simp5611_0[0:0], fa3_32min_0[0:0], fa3_32min_0[3:3], fa3_32min_0[5:5]);
  INV I645 (simp5611_0[1:1], fa3_32min_0[6:6]);
  NAND2 I646 (termf_3[32:32], simp5611_0[0:0], simp5611_0[1:1]);
  NOR3 I647 (simp5621_0[0:0], fa3_32min_0[1:1], fa3_32min_0[2:2], fa3_32min_0[4:4]);
  INV I648 (simp5621_0[1:1], fa3_32min_0[7:7]);
  NAND2 I649 (termt_3[32:32], simp5621_0[0:0], simp5621_0[1:1]);
  AO222 I650 (ct3__0[32:32], termt_1[32:32], termt_2[32:32], termt_1[32:32], ct3__0[31:31], termt_2[32:32], ct3__0[31:31]);
  AO222 I651 (cf3__0[32:32], termf_1[32:32], termf_2[32:32], termf_1[32:32], cf3__0[31:31], termf_2[32:32], cf3__0[31:31]);
  BUFF I652 (o_0r0[0:0], termf_3[0:0]);
  BUFF I653 (o_0r0[1:1], termf_3[1:1]);
  BUFF I654 (o_0r0[2:2], termf_3[2:2]);
  BUFF I655 (o_0r0[3:3], termf_3[3:3]);
  BUFF I656 (o_0r0[4:4], termf_3[4:4]);
  BUFF I657 (o_0r0[5:5], termf_3[5:5]);
  BUFF I658 (o_0r0[6:6], termf_3[6:6]);
  BUFF I659 (o_0r0[7:7], termf_3[7:7]);
  BUFF I660 (o_0r0[8:8], termf_3[8:8]);
  BUFF I661 (o_0r0[9:9], termf_3[9:9]);
  BUFF I662 (o_0r0[10:10], termf_3[10:10]);
  BUFF I663 (o_0r0[11:11], termf_3[11:11]);
  BUFF I664 (o_0r0[12:12], termf_3[12:12]);
  BUFF I665 (o_0r0[13:13], termf_3[13:13]);
  BUFF I666 (o_0r0[14:14], termf_3[14:14]);
  BUFF I667 (o_0r0[15:15], termf_3[15:15]);
  BUFF I668 (o_0r0[16:16], termf_3[16:16]);
  BUFF I669 (o_0r0[17:17], termf_3[17:17]);
  BUFF I670 (o_0r0[18:18], termf_3[18:18]);
  BUFF I671 (o_0r0[19:19], termf_3[19:19]);
  BUFF I672 (o_0r0[20:20], termf_3[20:20]);
  BUFF I673 (o_0r0[21:21], termf_3[21:21]);
  BUFF I674 (o_0r0[22:22], termf_3[22:22]);
  BUFF I675 (o_0r0[23:23], termf_3[23:23]);
  BUFF I676 (o_0r0[24:24], termf_3[24:24]);
  BUFF I677 (o_0r0[25:25], termf_3[25:25]);
  BUFF I678 (o_0r0[26:26], termf_3[26:26]);
  BUFF I679 (o_0r0[27:27], termf_3[27:27]);
  BUFF I680 (o_0r0[28:28], termf_3[28:28]);
  BUFF I681 (o_0r0[29:29], termf_3[29:29]);
  BUFF I682 (o_0r0[30:30], termf_3[30:30]);
  BUFF I683 (o_0r0[31:31], termf_3[31:31]);
  BUFF I684 (o_0r1[0:0], termt_3[0:0]);
  BUFF I685 (o_0r1[1:1], termt_3[1:1]);
  BUFF I686 (o_0r1[2:2], termt_3[2:2]);
  BUFF I687 (o_0r1[3:3], termt_3[3:3]);
  BUFF I688 (o_0r1[4:4], termt_3[4:4]);
  BUFF I689 (o_0r1[5:5], termt_3[5:5]);
  BUFF I690 (o_0r1[6:6], termt_3[6:6]);
  BUFF I691 (o_0r1[7:7], termt_3[7:7]);
  BUFF I692 (o_0r1[8:8], termt_3[8:8]);
  BUFF I693 (o_0r1[9:9], termt_3[9:9]);
  BUFF I694 (o_0r1[10:10], termt_3[10:10]);
  BUFF I695 (o_0r1[11:11], termt_3[11:11]);
  BUFF I696 (o_0r1[12:12], termt_3[12:12]);
  BUFF I697 (o_0r1[13:13], termt_3[13:13]);
  BUFF I698 (o_0r1[14:14], termt_3[14:14]);
  BUFF I699 (o_0r1[15:15], termt_3[15:15]);
  BUFF I700 (o_0r1[16:16], termt_3[16:16]);
  BUFF I701 (o_0r1[17:17], termt_3[17:17]);
  BUFF I702 (o_0r1[18:18], termt_3[18:18]);
  BUFF I703 (o_0r1[19:19], termt_3[19:19]);
  BUFF I704 (o_0r1[20:20], termt_3[20:20]);
  BUFF I705 (o_0r1[21:21], termt_3[21:21]);
  BUFF I706 (o_0r1[22:22], termt_3[22:22]);
  BUFF I707 (o_0r1[23:23], termt_3[23:23]);
  BUFF I708 (o_0r1[24:24], termt_3[24:24]);
  BUFF I709 (o_0r1[25:25], termt_3[25:25]);
  BUFF I710 (o_0r1[26:26], termt_3[26:26]);
  BUFF I711 (o_0r1[27:27], termt_3[27:27]);
  BUFF I712 (o_0r1[28:28], termt_3[28:28]);
  BUFF I713 (o_0r1[29:29], termt_3[29:29]);
  BUFF I714 (o_0r1[30:30], termt_3[30:30]);
  BUFF I715 (o_0r1[31:31], termt_3[31:31]);
  BUFF I716 (i_0a, o_0a);
endmodule

// latch tkl32x1 width = 32, depth = 1
module tkl32x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [31:0] bcomp_0;
  wire [10:0] simp991_0;
  wire [3:0] simp992_0;
  wire [1:0] simp993_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r0[10:10], i_0r0[10:10], bna_0, reset);
  C2R I11 (o_0r0[11:11], i_0r0[11:11], bna_0, reset);
  C2R I12 (o_0r0[12:12], i_0r0[12:12], bna_0, reset);
  C2R I13 (o_0r0[13:13], i_0r0[13:13], bna_0, reset);
  C2R I14 (o_0r0[14:14], i_0r0[14:14], bna_0, reset);
  C2R I15 (o_0r0[15:15], i_0r0[15:15], bna_0, reset);
  C2R I16 (o_0r0[16:16], i_0r0[16:16], bna_0, reset);
  C2R I17 (o_0r0[17:17], i_0r0[17:17], bna_0, reset);
  C2R I18 (o_0r0[18:18], i_0r0[18:18], bna_0, reset);
  C2R I19 (o_0r0[19:19], i_0r0[19:19], bna_0, reset);
  C2R I20 (o_0r0[20:20], i_0r0[20:20], bna_0, reset);
  C2R I21 (o_0r0[21:21], i_0r0[21:21], bna_0, reset);
  C2R I22 (o_0r0[22:22], i_0r0[22:22], bna_0, reset);
  C2R I23 (o_0r0[23:23], i_0r0[23:23], bna_0, reset);
  C2R I24 (o_0r0[24:24], i_0r0[24:24], bna_0, reset);
  C2R I25 (o_0r0[25:25], i_0r0[25:25], bna_0, reset);
  C2R I26 (o_0r0[26:26], i_0r0[26:26], bna_0, reset);
  C2R I27 (o_0r0[27:27], i_0r0[27:27], bna_0, reset);
  C2R I28 (o_0r0[28:28], i_0r0[28:28], bna_0, reset);
  C2R I29 (o_0r0[29:29], i_0r0[29:29], bna_0, reset);
  C2R I30 (o_0r0[30:30], i_0r0[30:30], bna_0, reset);
  C2R I31 (o_0r0[31:31], i_0r0[31:31], bna_0, reset);
  C2R I32 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I33 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I34 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I35 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I36 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I37 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I38 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I39 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I40 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I41 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  C2R I42 (o_0r1[10:10], i_0r1[10:10], bna_0, reset);
  C2R I43 (o_0r1[11:11], i_0r1[11:11], bna_0, reset);
  C2R I44 (o_0r1[12:12], i_0r1[12:12], bna_0, reset);
  C2R I45 (o_0r1[13:13], i_0r1[13:13], bna_0, reset);
  C2R I46 (o_0r1[14:14], i_0r1[14:14], bna_0, reset);
  C2R I47 (o_0r1[15:15], i_0r1[15:15], bna_0, reset);
  C2R I48 (o_0r1[16:16], i_0r1[16:16], bna_0, reset);
  C2R I49 (o_0r1[17:17], i_0r1[17:17], bna_0, reset);
  C2R I50 (o_0r1[18:18], i_0r1[18:18], bna_0, reset);
  C2R I51 (o_0r1[19:19], i_0r1[19:19], bna_0, reset);
  C2R I52 (o_0r1[20:20], i_0r1[20:20], bna_0, reset);
  C2R I53 (o_0r1[21:21], i_0r1[21:21], bna_0, reset);
  C2R I54 (o_0r1[22:22], i_0r1[22:22], bna_0, reset);
  C2R I55 (o_0r1[23:23], i_0r1[23:23], bna_0, reset);
  C2R I56 (o_0r1[24:24], i_0r1[24:24], bna_0, reset);
  C2R I57 (o_0r1[25:25], i_0r1[25:25], bna_0, reset);
  C2R I58 (o_0r1[26:26], i_0r1[26:26], bna_0, reset);
  C2R I59 (o_0r1[27:27], i_0r1[27:27], bna_0, reset);
  C2R I60 (o_0r1[28:28], i_0r1[28:28], bna_0, reset);
  C2R I61 (o_0r1[29:29], i_0r1[29:29], bna_0, reset);
  C2R I62 (o_0r1[30:30], i_0r1[30:30], bna_0, reset);
  C2R I63 (o_0r1[31:31], i_0r1[31:31], bna_0, reset);
  INV I64 (bna_0, o_0a);
  OR2 I65 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I66 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I67 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I68 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I69 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I70 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I71 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I72 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I73 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I74 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  OR2 I75 (bcomp_0[10:10], o_0r0[10:10], o_0r1[10:10]);
  OR2 I76 (bcomp_0[11:11], o_0r0[11:11], o_0r1[11:11]);
  OR2 I77 (bcomp_0[12:12], o_0r0[12:12], o_0r1[12:12]);
  OR2 I78 (bcomp_0[13:13], o_0r0[13:13], o_0r1[13:13]);
  OR2 I79 (bcomp_0[14:14], o_0r0[14:14], o_0r1[14:14]);
  OR2 I80 (bcomp_0[15:15], o_0r0[15:15], o_0r1[15:15]);
  OR2 I81 (bcomp_0[16:16], o_0r0[16:16], o_0r1[16:16]);
  OR2 I82 (bcomp_0[17:17], o_0r0[17:17], o_0r1[17:17]);
  OR2 I83 (bcomp_0[18:18], o_0r0[18:18], o_0r1[18:18]);
  OR2 I84 (bcomp_0[19:19], o_0r0[19:19], o_0r1[19:19]);
  OR2 I85 (bcomp_0[20:20], o_0r0[20:20], o_0r1[20:20]);
  OR2 I86 (bcomp_0[21:21], o_0r0[21:21], o_0r1[21:21]);
  OR2 I87 (bcomp_0[22:22], o_0r0[22:22], o_0r1[22:22]);
  OR2 I88 (bcomp_0[23:23], o_0r0[23:23], o_0r1[23:23]);
  OR2 I89 (bcomp_0[24:24], o_0r0[24:24], o_0r1[24:24]);
  OR2 I90 (bcomp_0[25:25], o_0r0[25:25], o_0r1[25:25]);
  OR2 I91 (bcomp_0[26:26], o_0r0[26:26], o_0r1[26:26]);
  OR2 I92 (bcomp_0[27:27], o_0r0[27:27], o_0r1[27:27]);
  OR2 I93 (bcomp_0[28:28], o_0r0[28:28], o_0r1[28:28]);
  OR2 I94 (bcomp_0[29:29], o_0r0[29:29], o_0r1[29:29]);
  OR2 I95 (bcomp_0[30:30], o_0r0[30:30], o_0r1[30:30]);
  OR2 I96 (bcomp_0[31:31], o_0r0[31:31], o_0r1[31:31]);
  C3 I97 (simp991_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I98 (simp991_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I99 (simp991_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  C3 I100 (simp991_0[3:3], bcomp_0[9:9], bcomp_0[10:10], bcomp_0[11:11]);
  C3 I101 (simp991_0[4:4], bcomp_0[12:12], bcomp_0[13:13], bcomp_0[14:14]);
  C3 I102 (simp991_0[5:5], bcomp_0[15:15], bcomp_0[16:16], bcomp_0[17:17]);
  C3 I103 (simp991_0[6:6], bcomp_0[18:18], bcomp_0[19:19], bcomp_0[20:20]);
  C3 I104 (simp991_0[7:7], bcomp_0[21:21], bcomp_0[22:22], bcomp_0[23:23]);
  C3 I105 (simp991_0[8:8], bcomp_0[24:24], bcomp_0[25:25], bcomp_0[26:26]);
  C3 I106 (simp991_0[9:9], bcomp_0[27:27], bcomp_0[28:28], bcomp_0[29:29]);
  C2 I107 (simp991_0[10:10], bcomp_0[30:30], bcomp_0[31:31]);
  C3 I108 (simp992_0[0:0], simp991_0[0:0], simp991_0[1:1], simp991_0[2:2]);
  C3 I109 (simp992_0[1:1], simp991_0[3:3], simp991_0[4:4], simp991_0[5:5]);
  C3 I110 (simp992_0[2:2], simp991_0[6:6], simp991_0[7:7], simp991_0[8:8]);
  C2 I111 (simp992_0[3:3], simp991_0[9:9], simp991_0[10:10]);
  C3 I112 (simp993_0[0:0], simp992_0[0:0], simp992_0[1:1], simp992_0[2:2]);
  BUFF I113 (simp993_0[1:1], simp992_0[3:3]);
  C2 I114 (i_0a, simp993_0[0:0], simp993_0[1:1]);
endmodule

// latch tkl0x1 width = 0, depth = 1
module tkl0x1 (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire b_0;
  C2R I0 (o_0r, i_0r, b_0, reset);
  INV I1 (b_0, o_0a);
  BUFF I2 (i_0a, o_0r);
endmodule

// latch tkl4x1 width = 4, depth = 1
module tkl4x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [3:0] bcomp_0;
  wire [1:0] simp151_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I5 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I6 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I7 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  INV I8 (bna_0, o_0a);
  OR2 I9 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I10 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I11 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I12 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  C3 I13 (simp151_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  BUFF I14 (simp151_0[1:1], bcomp_0[3:3]);
  C2 I15 (i_0a, simp151_0[0:0], simp151_0[1:1]);
endmodule

// latch tkl64x1 width = 64, depth = 1
module tkl64x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [63:0] o_0r0;
  output [63:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [63:0] bcomp_0;
  wire [21:0] simp1951_0;
  wire [7:0] simp1952_0;
  wire [2:0] simp1953_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r0[10:10], i_0r0[10:10], bna_0, reset);
  C2R I11 (o_0r0[11:11], i_0r0[11:11], bna_0, reset);
  C2R I12 (o_0r0[12:12], i_0r0[12:12], bna_0, reset);
  C2R I13 (o_0r0[13:13], i_0r0[13:13], bna_0, reset);
  C2R I14 (o_0r0[14:14], i_0r0[14:14], bna_0, reset);
  C2R I15 (o_0r0[15:15], i_0r0[15:15], bna_0, reset);
  C2R I16 (o_0r0[16:16], i_0r0[16:16], bna_0, reset);
  C2R I17 (o_0r0[17:17], i_0r0[17:17], bna_0, reset);
  C2R I18 (o_0r0[18:18], i_0r0[18:18], bna_0, reset);
  C2R I19 (o_0r0[19:19], i_0r0[19:19], bna_0, reset);
  C2R I20 (o_0r0[20:20], i_0r0[20:20], bna_0, reset);
  C2R I21 (o_0r0[21:21], i_0r0[21:21], bna_0, reset);
  C2R I22 (o_0r0[22:22], i_0r0[22:22], bna_0, reset);
  C2R I23 (o_0r0[23:23], i_0r0[23:23], bna_0, reset);
  C2R I24 (o_0r0[24:24], i_0r0[24:24], bna_0, reset);
  C2R I25 (o_0r0[25:25], i_0r0[25:25], bna_0, reset);
  C2R I26 (o_0r0[26:26], i_0r0[26:26], bna_0, reset);
  C2R I27 (o_0r0[27:27], i_0r0[27:27], bna_0, reset);
  C2R I28 (o_0r0[28:28], i_0r0[28:28], bna_0, reset);
  C2R I29 (o_0r0[29:29], i_0r0[29:29], bna_0, reset);
  C2R I30 (o_0r0[30:30], i_0r0[30:30], bna_0, reset);
  C2R I31 (o_0r0[31:31], i_0r0[31:31], bna_0, reset);
  C2R I32 (o_0r0[32:32], i_0r0[32:32], bna_0, reset);
  C2R I33 (o_0r0[33:33], i_0r0[33:33], bna_0, reset);
  C2R I34 (o_0r0[34:34], i_0r0[34:34], bna_0, reset);
  C2R I35 (o_0r0[35:35], i_0r0[35:35], bna_0, reset);
  C2R I36 (o_0r0[36:36], i_0r0[36:36], bna_0, reset);
  C2R I37 (o_0r0[37:37], i_0r0[37:37], bna_0, reset);
  C2R I38 (o_0r0[38:38], i_0r0[38:38], bna_0, reset);
  C2R I39 (o_0r0[39:39], i_0r0[39:39], bna_0, reset);
  C2R I40 (o_0r0[40:40], i_0r0[40:40], bna_0, reset);
  C2R I41 (o_0r0[41:41], i_0r0[41:41], bna_0, reset);
  C2R I42 (o_0r0[42:42], i_0r0[42:42], bna_0, reset);
  C2R I43 (o_0r0[43:43], i_0r0[43:43], bna_0, reset);
  C2R I44 (o_0r0[44:44], i_0r0[44:44], bna_0, reset);
  C2R I45 (o_0r0[45:45], i_0r0[45:45], bna_0, reset);
  C2R I46 (o_0r0[46:46], i_0r0[46:46], bna_0, reset);
  C2R I47 (o_0r0[47:47], i_0r0[47:47], bna_0, reset);
  C2R I48 (o_0r0[48:48], i_0r0[48:48], bna_0, reset);
  C2R I49 (o_0r0[49:49], i_0r0[49:49], bna_0, reset);
  C2R I50 (o_0r0[50:50], i_0r0[50:50], bna_0, reset);
  C2R I51 (o_0r0[51:51], i_0r0[51:51], bna_0, reset);
  C2R I52 (o_0r0[52:52], i_0r0[52:52], bna_0, reset);
  C2R I53 (o_0r0[53:53], i_0r0[53:53], bna_0, reset);
  C2R I54 (o_0r0[54:54], i_0r0[54:54], bna_0, reset);
  C2R I55 (o_0r0[55:55], i_0r0[55:55], bna_0, reset);
  C2R I56 (o_0r0[56:56], i_0r0[56:56], bna_0, reset);
  C2R I57 (o_0r0[57:57], i_0r0[57:57], bna_0, reset);
  C2R I58 (o_0r0[58:58], i_0r0[58:58], bna_0, reset);
  C2R I59 (o_0r0[59:59], i_0r0[59:59], bna_0, reset);
  C2R I60 (o_0r0[60:60], i_0r0[60:60], bna_0, reset);
  C2R I61 (o_0r0[61:61], i_0r0[61:61], bna_0, reset);
  C2R I62 (o_0r0[62:62], i_0r0[62:62], bna_0, reset);
  C2R I63 (o_0r0[63:63], i_0r0[63:63], bna_0, reset);
  C2R I64 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I65 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I66 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I67 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I68 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I69 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I70 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I71 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I72 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I73 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  C2R I74 (o_0r1[10:10], i_0r1[10:10], bna_0, reset);
  C2R I75 (o_0r1[11:11], i_0r1[11:11], bna_0, reset);
  C2R I76 (o_0r1[12:12], i_0r1[12:12], bna_0, reset);
  C2R I77 (o_0r1[13:13], i_0r1[13:13], bna_0, reset);
  C2R I78 (o_0r1[14:14], i_0r1[14:14], bna_0, reset);
  C2R I79 (o_0r1[15:15], i_0r1[15:15], bna_0, reset);
  C2R I80 (o_0r1[16:16], i_0r1[16:16], bna_0, reset);
  C2R I81 (o_0r1[17:17], i_0r1[17:17], bna_0, reset);
  C2R I82 (o_0r1[18:18], i_0r1[18:18], bna_0, reset);
  C2R I83 (o_0r1[19:19], i_0r1[19:19], bna_0, reset);
  C2R I84 (o_0r1[20:20], i_0r1[20:20], bna_0, reset);
  C2R I85 (o_0r1[21:21], i_0r1[21:21], bna_0, reset);
  C2R I86 (o_0r1[22:22], i_0r1[22:22], bna_0, reset);
  C2R I87 (o_0r1[23:23], i_0r1[23:23], bna_0, reset);
  C2R I88 (o_0r1[24:24], i_0r1[24:24], bna_0, reset);
  C2R I89 (o_0r1[25:25], i_0r1[25:25], bna_0, reset);
  C2R I90 (o_0r1[26:26], i_0r1[26:26], bna_0, reset);
  C2R I91 (o_0r1[27:27], i_0r1[27:27], bna_0, reset);
  C2R I92 (o_0r1[28:28], i_0r1[28:28], bna_0, reset);
  C2R I93 (o_0r1[29:29], i_0r1[29:29], bna_0, reset);
  C2R I94 (o_0r1[30:30], i_0r1[30:30], bna_0, reset);
  C2R I95 (o_0r1[31:31], i_0r1[31:31], bna_0, reset);
  C2R I96 (o_0r1[32:32], i_0r1[32:32], bna_0, reset);
  C2R I97 (o_0r1[33:33], i_0r1[33:33], bna_0, reset);
  C2R I98 (o_0r1[34:34], i_0r1[34:34], bna_0, reset);
  C2R I99 (o_0r1[35:35], i_0r1[35:35], bna_0, reset);
  C2R I100 (o_0r1[36:36], i_0r1[36:36], bna_0, reset);
  C2R I101 (o_0r1[37:37], i_0r1[37:37], bna_0, reset);
  C2R I102 (o_0r1[38:38], i_0r1[38:38], bna_0, reset);
  C2R I103 (o_0r1[39:39], i_0r1[39:39], bna_0, reset);
  C2R I104 (o_0r1[40:40], i_0r1[40:40], bna_0, reset);
  C2R I105 (o_0r1[41:41], i_0r1[41:41], bna_0, reset);
  C2R I106 (o_0r1[42:42], i_0r1[42:42], bna_0, reset);
  C2R I107 (o_0r1[43:43], i_0r1[43:43], bna_0, reset);
  C2R I108 (o_0r1[44:44], i_0r1[44:44], bna_0, reset);
  C2R I109 (o_0r1[45:45], i_0r1[45:45], bna_0, reset);
  C2R I110 (o_0r1[46:46], i_0r1[46:46], bna_0, reset);
  C2R I111 (o_0r1[47:47], i_0r1[47:47], bna_0, reset);
  C2R I112 (o_0r1[48:48], i_0r1[48:48], bna_0, reset);
  C2R I113 (o_0r1[49:49], i_0r1[49:49], bna_0, reset);
  C2R I114 (o_0r1[50:50], i_0r1[50:50], bna_0, reset);
  C2R I115 (o_0r1[51:51], i_0r1[51:51], bna_0, reset);
  C2R I116 (o_0r1[52:52], i_0r1[52:52], bna_0, reset);
  C2R I117 (o_0r1[53:53], i_0r1[53:53], bna_0, reset);
  C2R I118 (o_0r1[54:54], i_0r1[54:54], bna_0, reset);
  C2R I119 (o_0r1[55:55], i_0r1[55:55], bna_0, reset);
  C2R I120 (o_0r1[56:56], i_0r1[56:56], bna_0, reset);
  C2R I121 (o_0r1[57:57], i_0r1[57:57], bna_0, reset);
  C2R I122 (o_0r1[58:58], i_0r1[58:58], bna_0, reset);
  C2R I123 (o_0r1[59:59], i_0r1[59:59], bna_0, reset);
  C2R I124 (o_0r1[60:60], i_0r1[60:60], bna_0, reset);
  C2R I125 (o_0r1[61:61], i_0r1[61:61], bna_0, reset);
  C2R I126 (o_0r1[62:62], i_0r1[62:62], bna_0, reset);
  C2R I127 (o_0r1[63:63], i_0r1[63:63], bna_0, reset);
  INV I128 (bna_0, o_0a);
  OR2 I129 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I130 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I131 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I132 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I133 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I134 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I135 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I136 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I137 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I138 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  OR2 I139 (bcomp_0[10:10], o_0r0[10:10], o_0r1[10:10]);
  OR2 I140 (bcomp_0[11:11], o_0r0[11:11], o_0r1[11:11]);
  OR2 I141 (bcomp_0[12:12], o_0r0[12:12], o_0r1[12:12]);
  OR2 I142 (bcomp_0[13:13], o_0r0[13:13], o_0r1[13:13]);
  OR2 I143 (bcomp_0[14:14], o_0r0[14:14], o_0r1[14:14]);
  OR2 I144 (bcomp_0[15:15], o_0r0[15:15], o_0r1[15:15]);
  OR2 I145 (bcomp_0[16:16], o_0r0[16:16], o_0r1[16:16]);
  OR2 I146 (bcomp_0[17:17], o_0r0[17:17], o_0r1[17:17]);
  OR2 I147 (bcomp_0[18:18], o_0r0[18:18], o_0r1[18:18]);
  OR2 I148 (bcomp_0[19:19], o_0r0[19:19], o_0r1[19:19]);
  OR2 I149 (bcomp_0[20:20], o_0r0[20:20], o_0r1[20:20]);
  OR2 I150 (bcomp_0[21:21], o_0r0[21:21], o_0r1[21:21]);
  OR2 I151 (bcomp_0[22:22], o_0r0[22:22], o_0r1[22:22]);
  OR2 I152 (bcomp_0[23:23], o_0r0[23:23], o_0r1[23:23]);
  OR2 I153 (bcomp_0[24:24], o_0r0[24:24], o_0r1[24:24]);
  OR2 I154 (bcomp_0[25:25], o_0r0[25:25], o_0r1[25:25]);
  OR2 I155 (bcomp_0[26:26], o_0r0[26:26], o_0r1[26:26]);
  OR2 I156 (bcomp_0[27:27], o_0r0[27:27], o_0r1[27:27]);
  OR2 I157 (bcomp_0[28:28], o_0r0[28:28], o_0r1[28:28]);
  OR2 I158 (bcomp_0[29:29], o_0r0[29:29], o_0r1[29:29]);
  OR2 I159 (bcomp_0[30:30], o_0r0[30:30], o_0r1[30:30]);
  OR2 I160 (bcomp_0[31:31], o_0r0[31:31], o_0r1[31:31]);
  OR2 I161 (bcomp_0[32:32], o_0r0[32:32], o_0r1[32:32]);
  OR2 I162 (bcomp_0[33:33], o_0r0[33:33], o_0r1[33:33]);
  OR2 I163 (bcomp_0[34:34], o_0r0[34:34], o_0r1[34:34]);
  OR2 I164 (bcomp_0[35:35], o_0r0[35:35], o_0r1[35:35]);
  OR2 I165 (bcomp_0[36:36], o_0r0[36:36], o_0r1[36:36]);
  OR2 I166 (bcomp_0[37:37], o_0r0[37:37], o_0r1[37:37]);
  OR2 I167 (bcomp_0[38:38], o_0r0[38:38], o_0r1[38:38]);
  OR2 I168 (bcomp_0[39:39], o_0r0[39:39], o_0r1[39:39]);
  OR2 I169 (bcomp_0[40:40], o_0r0[40:40], o_0r1[40:40]);
  OR2 I170 (bcomp_0[41:41], o_0r0[41:41], o_0r1[41:41]);
  OR2 I171 (bcomp_0[42:42], o_0r0[42:42], o_0r1[42:42]);
  OR2 I172 (bcomp_0[43:43], o_0r0[43:43], o_0r1[43:43]);
  OR2 I173 (bcomp_0[44:44], o_0r0[44:44], o_0r1[44:44]);
  OR2 I174 (bcomp_0[45:45], o_0r0[45:45], o_0r1[45:45]);
  OR2 I175 (bcomp_0[46:46], o_0r0[46:46], o_0r1[46:46]);
  OR2 I176 (bcomp_0[47:47], o_0r0[47:47], o_0r1[47:47]);
  OR2 I177 (bcomp_0[48:48], o_0r0[48:48], o_0r1[48:48]);
  OR2 I178 (bcomp_0[49:49], o_0r0[49:49], o_0r1[49:49]);
  OR2 I179 (bcomp_0[50:50], o_0r0[50:50], o_0r1[50:50]);
  OR2 I180 (bcomp_0[51:51], o_0r0[51:51], o_0r1[51:51]);
  OR2 I181 (bcomp_0[52:52], o_0r0[52:52], o_0r1[52:52]);
  OR2 I182 (bcomp_0[53:53], o_0r0[53:53], o_0r1[53:53]);
  OR2 I183 (bcomp_0[54:54], o_0r0[54:54], o_0r1[54:54]);
  OR2 I184 (bcomp_0[55:55], o_0r0[55:55], o_0r1[55:55]);
  OR2 I185 (bcomp_0[56:56], o_0r0[56:56], o_0r1[56:56]);
  OR2 I186 (bcomp_0[57:57], o_0r0[57:57], o_0r1[57:57]);
  OR2 I187 (bcomp_0[58:58], o_0r0[58:58], o_0r1[58:58]);
  OR2 I188 (bcomp_0[59:59], o_0r0[59:59], o_0r1[59:59]);
  OR2 I189 (bcomp_0[60:60], o_0r0[60:60], o_0r1[60:60]);
  OR2 I190 (bcomp_0[61:61], o_0r0[61:61], o_0r1[61:61]);
  OR2 I191 (bcomp_0[62:62], o_0r0[62:62], o_0r1[62:62]);
  OR2 I192 (bcomp_0[63:63], o_0r0[63:63], o_0r1[63:63]);
  C3 I193 (simp1951_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I194 (simp1951_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I195 (simp1951_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  C3 I196 (simp1951_0[3:3], bcomp_0[9:9], bcomp_0[10:10], bcomp_0[11:11]);
  C3 I197 (simp1951_0[4:4], bcomp_0[12:12], bcomp_0[13:13], bcomp_0[14:14]);
  C3 I198 (simp1951_0[5:5], bcomp_0[15:15], bcomp_0[16:16], bcomp_0[17:17]);
  C3 I199 (simp1951_0[6:6], bcomp_0[18:18], bcomp_0[19:19], bcomp_0[20:20]);
  C3 I200 (simp1951_0[7:7], bcomp_0[21:21], bcomp_0[22:22], bcomp_0[23:23]);
  C3 I201 (simp1951_0[8:8], bcomp_0[24:24], bcomp_0[25:25], bcomp_0[26:26]);
  C3 I202 (simp1951_0[9:9], bcomp_0[27:27], bcomp_0[28:28], bcomp_0[29:29]);
  C3 I203 (simp1951_0[10:10], bcomp_0[30:30], bcomp_0[31:31], bcomp_0[32:32]);
  C3 I204 (simp1951_0[11:11], bcomp_0[33:33], bcomp_0[34:34], bcomp_0[35:35]);
  C3 I205 (simp1951_0[12:12], bcomp_0[36:36], bcomp_0[37:37], bcomp_0[38:38]);
  C3 I206 (simp1951_0[13:13], bcomp_0[39:39], bcomp_0[40:40], bcomp_0[41:41]);
  C3 I207 (simp1951_0[14:14], bcomp_0[42:42], bcomp_0[43:43], bcomp_0[44:44]);
  C3 I208 (simp1951_0[15:15], bcomp_0[45:45], bcomp_0[46:46], bcomp_0[47:47]);
  C3 I209 (simp1951_0[16:16], bcomp_0[48:48], bcomp_0[49:49], bcomp_0[50:50]);
  C3 I210 (simp1951_0[17:17], bcomp_0[51:51], bcomp_0[52:52], bcomp_0[53:53]);
  C3 I211 (simp1951_0[18:18], bcomp_0[54:54], bcomp_0[55:55], bcomp_0[56:56]);
  C3 I212 (simp1951_0[19:19], bcomp_0[57:57], bcomp_0[58:58], bcomp_0[59:59]);
  C3 I213 (simp1951_0[20:20], bcomp_0[60:60], bcomp_0[61:61], bcomp_0[62:62]);
  BUFF I214 (simp1951_0[21:21], bcomp_0[63:63]);
  C3 I215 (simp1952_0[0:0], simp1951_0[0:0], simp1951_0[1:1], simp1951_0[2:2]);
  C3 I216 (simp1952_0[1:1], simp1951_0[3:3], simp1951_0[4:4], simp1951_0[5:5]);
  C3 I217 (simp1952_0[2:2], simp1951_0[6:6], simp1951_0[7:7], simp1951_0[8:8]);
  C3 I218 (simp1952_0[3:3], simp1951_0[9:9], simp1951_0[10:10], simp1951_0[11:11]);
  C3 I219 (simp1952_0[4:4], simp1951_0[12:12], simp1951_0[13:13], simp1951_0[14:14]);
  C3 I220 (simp1952_0[5:5], simp1951_0[15:15], simp1951_0[16:16], simp1951_0[17:17]);
  C3 I221 (simp1952_0[6:6], simp1951_0[18:18], simp1951_0[19:19], simp1951_0[20:20]);
  BUFF I222 (simp1952_0[7:7], simp1951_0[21:21]);
  C3 I223 (simp1953_0[0:0], simp1952_0[0:0], simp1952_0[1:1], simp1952_0[2:2]);
  C3 I224 (simp1953_0[1:1], simp1952_0[3:3], simp1952_0[4:4], simp1952_0[5:5]);
  C2 I225 (simp1953_0[2:2], simp1952_0[6:6], simp1952_0[7:7]);
  C3 I226 (i_0a, simp1953_0[0:0], simp1953_0[1:1], simp1953_0[2:2]);
endmodule

// latch tkl33x1 width = 33, depth = 1
module tkl33x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [32:0] bcomp_0;
  wire [10:0] simp1021_0;
  wire [3:0] simp1022_0;
  wire [1:0] simp1023_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r0[10:10], i_0r0[10:10], bna_0, reset);
  C2R I11 (o_0r0[11:11], i_0r0[11:11], bna_0, reset);
  C2R I12 (o_0r0[12:12], i_0r0[12:12], bna_0, reset);
  C2R I13 (o_0r0[13:13], i_0r0[13:13], bna_0, reset);
  C2R I14 (o_0r0[14:14], i_0r0[14:14], bna_0, reset);
  C2R I15 (o_0r0[15:15], i_0r0[15:15], bna_0, reset);
  C2R I16 (o_0r0[16:16], i_0r0[16:16], bna_0, reset);
  C2R I17 (o_0r0[17:17], i_0r0[17:17], bna_0, reset);
  C2R I18 (o_0r0[18:18], i_0r0[18:18], bna_0, reset);
  C2R I19 (o_0r0[19:19], i_0r0[19:19], bna_0, reset);
  C2R I20 (o_0r0[20:20], i_0r0[20:20], bna_0, reset);
  C2R I21 (o_0r0[21:21], i_0r0[21:21], bna_0, reset);
  C2R I22 (o_0r0[22:22], i_0r0[22:22], bna_0, reset);
  C2R I23 (o_0r0[23:23], i_0r0[23:23], bna_0, reset);
  C2R I24 (o_0r0[24:24], i_0r0[24:24], bna_0, reset);
  C2R I25 (o_0r0[25:25], i_0r0[25:25], bna_0, reset);
  C2R I26 (o_0r0[26:26], i_0r0[26:26], bna_0, reset);
  C2R I27 (o_0r0[27:27], i_0r0[27:27], bna_0, reset);
  C2R I28 (o_0r0[28:28], i_0r0[28:28], bna_0, reset);
  C2R I29 (o_0r0[29:29], i_0r0[29:29], bna_0, reset);
  C2R I30 (o_0r0[30:30], i_0r0[30:30], bna_0, reset);
  C2R I31 (o_0r0[31:31], i_0r0[31:31], bna_0, reset);
  C2R I32 (o_0r0[32:32], i_0r0[32:32], bna_0, reset);
  C2R I33 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I34 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I35 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I36 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I37 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I38 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I39 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I40 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I41 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I42 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  C2R I43 (o_0r1[10:10], i_0r1[10:10], bna_0, reset);
  C2R I44 (o_0r1[11:11], i_0r1[11:11], bna_0, reset);
  C2R I45 (o_0r1[12:12], i_0r1[12:12], bna_0, reset);
  C2R I46 (o_0r1[13:13], i_0r1[13:13], bna_0, reset);
  C2R I47 (o_0r1[14:14], i_0r1[14:14], bna_0, reset);
  C2R I48 (o_0r1[15:15], i_0r1[15:15], bna_0, reset);
  C2R I49 (o_0r1[16:16], i_0r1[16:16], bna_0, reset);
  C2R I50 (o_0r1[17:17], i_0r1[17:17], bna_0, reset);
  C2R I51 (o_0r1[18:18], i_0r1[18:18], bna_0, reset);
  C2R I52 (o_0r1[19:19], i_0r1[19:19], bna_0, reset);
  C2R I53 (o_0r1[20:20], i_0r1[20:20], bna_0, reset);
  C2R I54 (o_0r1[21:21], i_0r1[21:21], bna_0, reset);
  C2R I55 (o_0r1[22:22], i_0r1[22:22], bna_0, reset);
  C2R I56 (o_0r1[23:23], i_0r1[23:23], bna_0, reset);
  C2R I57 (o_0r1[24:24], i_0r1[24:24], bna_0, reset);
  C2R I58 (o_0r1[25:25], i_0r1[25:25], bna_0, reset);
  C2R I59 (o_0r1[26:26], i_0r1[26:26], bna_0, reset);
  C2R I60 (o_0r1[27:27], i_0r1[27:27], bna_0, reset);
  C2R I61 (o_0r1[28:28], i_0r1[28:28], bna_0, reset);
  C2R I62 (o_0r1[29:29], i_0r1[29:29], bna_0, reset);
  C2R I63 (o_0r1[30:30], i_0r1[30:30], bna_0, reset);
  C2R I64 (o_0r1[31:31], i_0r1[31:31], bna_0, reset);
  C2R I65 (o_0r1[32:32], i_0r1[32:32], bna_0, reset);
  INV I66 (bna_0, o_0a);
  OR2 I67 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I68 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I69 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I70 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I71 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I72 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I73 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I74 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I75 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I76 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  OR2 I77 (bcomp_0[10:10], o_0r0[10:10], o_0r1[10:10]);
  OR2 I78 (bcomp_0[11:11], o_0r0[11:11], o_0r1[11:11]);
  OR2 I79 (bcomp_0[12:12], o_0r0[12:12], o_0r1[12:12]);
  OR2 I80 (bcomp_0[13:13], o_0r0[13:13], o_0r1[13:13]);
  OR2 I81 (bcomp_0[14:14], o_0r0[14:14], o_0r1[14:14]);
  OR2 I82 (bcomp_0[15:15], o_0r0[15:15], o_0r1[15:15]);
  OR2 I83 (bcomp_0[16:16], o_0r0[16:16], o_0r1[16:16]);
  OR2 I84 (bcomp_0[17:17], o_0r0[17:17], o_0r1[17:17]);
  OR2 I85 (bcomp_0[18:18], o_0r0[18:18], o_0r1[18:18]);
  OR2 I86 (bcomp_0[19:19], o_0r0[19:19], o_0r1[19:19]);
  OR2 I87 (bcomp_0[20:20], o_0r0[20:20], o_0r1[20:20]);
  OR2 I88 (bcomp_0[21:21], o_0r0[21:21], o_0r1[21:21]);
  OR2 I89 (bcomp_0[22:22], o_0r0[22:22], o_0r1[22:22]);
  OR2 I90 (bcomp_0[23:23], o_0r0[23:23], o_0r1[23:23]);
  OR2 I91 (bcomp_0[24:24], o_0r0[24:24], o_0r1[24:24]);
  OR2 I92 (bcomp_0[25:25], o_0r0[25:25], o_0r1[25:25]);
  OR2 I93 (bcomp_0[26:26], o_0r0[26:26], o_0r1[26:26]);
  OR2 I94 (bcomp_0[27:27], o_0r0[27:27], o_0r1[27:27]);
  OR2 I95 (bcomp_0[28:28], o_0r0[28:28], o_0r1[28:28]);
  OR2 I96 (bcomp_0[29:29], o_0r0[29:29], o_0r1[29:29]);
  OR2 I97 (bcomp_0[30:30], o_0r0[30:30], o_0r1[30:30]);
  OR2 I98 (bcomp_0[31:31], o_0r0[31:31], o_0r1[31:31]);
  OR2 I99 (bcomp_0[32:32], o_0r0[32:32], o_0r1[32:32]);
  C3 I100 (simp1021_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I101 (simp1021_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I102 (simp1021_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  C3 I103 (simp1021_0[3:3], bcomp_0[9:9], bcomp_0[10:10], bcomp_0[11:11]);
  C3 I104 (simp1021_0[4:4], bcomp_0[12:12], bcomp_0[13:13], bcomp_0[14:14]);
  C3 I105 (simp1021_0[5:5], bcomp_0[15:15], bcomp_0[16:16], bcomp_0[17:17]);
  C3 I106 (simp1021_0[6:6], bcomp_0[18:18], bcomp_0[19:19], bcomp_0[20:20]);
  C3 I107 (simp1021_0[7:7], bcomp_0[21:21], bcomp_0[22:22], bcomp_0[23:23]);
  C3 I108 (simp1021_0[8:8], bcomp_0[24:24], bcomp_0[25:25], bcomp_0[26:26]);
  C3 I109 (simp1021_0[9:9], bcomp_0[27:27], bcomp_0[28:28], bcomp_0[29:29]);
  C3 I110 (simp1021_0[10:10], bcomp_0[30:30], bcomp_0[31:31], bcomp_0[32:32]);
  C3 I111 (simp1022_0[0:0], simp1021_0[0:0], simp1021_0[1:1], simp1021_0[2:2]);
  C3 I112 (simp1022_0[1:1], simp1021_0[3:3], simp1021_0[4:4], simp1021_0[5:5]);
  C3 I113 (simp1022_0[2:2], simp1021_0[6:6], simp1021_0[7:7], simp1021_0[8:8]);
  C2 I114 (simp1022_0[3:3], simp1021_0[9:9], simp1021_0[10:10]);
  C3 I115 (simp1023_0[0:0], simp1022_0[0:0], simp1022_0[1:1], simp1022_0[2:2]);
  BUFF I116 (simp1023_0[1:1], simp1022_0[3:3]);
  C2 I117 (i_0a, simp1023_0[0:0], simp1023_0[1:1]);
endmodule

// latch tkl3x1 width = 3, depth = 1
module tkl3x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [2:0] bcomp_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I4 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I5 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  INV I6 (bna_0, o_0a);
  OR2 I7 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I8 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I9 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  C3 I10 (i_0a, bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
endmodule

// latch tkl2x1 width = 2, depth = 1
module tkl2x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [1:0] bcomp_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I3 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  INV I4 (bna_0, o_0a);
  OR2 I5 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I6 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  C2 I7 (i_0a, bcomp_0[0:0], bcomp_0[1:1]);
endmodule

// latch tkl1x1 width = 1, depth = 1
module tkl1x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire bcomp_0;
  C2R I0 (o_0r0, i_0r0, bna_0, reset);
  C2R I1 (o_0r1, i_0r1, bna_0, reset);
  INV I2 (bna_0, o_0a);
  OR2 I3 (bcomp_0, o_0r0, o_0r1);
  BUFF I4 (i_0a, bcomp_0);
endmodule

module teak_Poly_eval (x_0r0, x_0r1, x_0a, coefs_0_0r0, coefs_0_0r1, coefs_0_0a, coefs_1_0r0, coefs_1_0r1, coefs_1_0a, coefs_2_0r0, coefs_2_0r1, coefs_2_0a, a_0r0, a_0r1, a_0a, reset);
  input [31:0] x_0r0;
  input [31:0] x_0r1;
  output x_0a;
  input [31:0] coefs_0_0r0;
  input [31:0] coefs_0_0r1;
  output coefs_0_0a;
  input [31:0] coefs_1_0r0;
  input [31:0] coefs_1_0r1;
  output coefs_1_0a;
  input [31:0] coefs_2_0r0;
  input [31:0] coefs_2_0r1;
  output coefs_2_0a;
  output [31:0] a_0r0;
  output [31:0] a_0r1;
  input a_0a;
  input reset;
  wire [31:0] L4P_0r0;
  wire [31:0] L4P_0r1;
  wire L4P_0a;
  wire [31:0] L4A_0r0;
  wire [31:0] L4A_0r1;
  wire L4A_0a;
  wire L7_0r;
  wire L7_0a;
  wire [31:0] L8_0r0;
  wire [31:0] L8_0r1;
  wire L8_0a;
  wire L9_0r;
  wire L9_0a;
  wire L13P_0r;
  wire L13P_0a;
  wire L13A_0r;
  wire L13A_0a;
  wire L14P_0r;
  wire L14P_0a;
  wire L14A_0r;
  wire L14A_0a;
  wire L16P_0r;
  wire L16P_0a;
  wire L16A_0r;
  wire L16A_0a;
  wire L21_0r0;
  wire L21_0r1;
  wire L21_0a;
  wire L38_0r;
  wire L38_0a;
  wire [31:0] L39_0r0;
  wire [31:0] L39_0r1;
  wire L39_0a;
  wire L41_0r;
  wire L41_0a;
  wire L45_0r;
  wire L45_0a;
  wire L49P_0r;
  wire L49P_0a;
  wire L49A_0r;
  wire L49A_0a;
  wire L54_0r0;
  wire L54_0r1;
  wire L54_0a;
  wire L56P_0r;
  wire L56P_0a;
  wire L56A_0r;
  wire L56A_0a;
  wire L61_0r;
  wire L61_0a;
  wire L63P_0r;
  wire L63P_0a;
  wire L63A_0r;
  wire L63A_0a;
  wire [3:0] L68_0r0;
  wire [3:0] L68_0r1;
  wire L68_0a;
  wire L71_0r;
  wire L71_0a;
  wire L72P_0r;
  wire L72P_0a;
  wire L72A_0r;
  wire L72A_0a;
  wire L73P_0r;
  wire L73P_0a;
  wire L73A_0r;
  wire L73A_0a;
  wire L75P_0r;
  wire L75P_0a;
  wire L75A_0r;
  wire L75A_0a;
  wire L80_0r0;
  wire L80_0r1;
  wire L80_0a;
  wire L82P_0r;
  wire L82P_0a;
  wire L82A_0r;
  wire L82A_0a;
  wire L87_0r;
  wire L87_0a;
  wire L89P_0r;
  wire L89P_0a;
  wire L89A_0r;
  wire L89A_0a;
  wire [3:0] L94P_0r0;
  wire [3:0] L94P_0r1;
  wire L94P_0a;
  wire [3:0] L94A_0r0;
  wire [3:0] L94A_0r1;
  wire L94A_0a;
  wire L97_0r;
  wire L97_0a;
  wire L98P_0r;
  wire L98P_0a;
  wire L98A_0r;
  wire L98A_0a;
  wire L99P_0r;
  wire L99P_0a;
  wire L99A_0r;
  wire L99A_0a;
  wire L101P_0r;
  wire L101P_0a;
  wire L101A_0r;
  wire L101A_0a;
  wire L106_0r0;
  wire L106_0r1;
  wire L106_0a;
  wire L110P_0r;
  wire L110P_0a;
  wire L110A_0r;
  wire L110A_0a;
  wire [31:0] L111P_0r0;
  wire [31:0] L111P_0r1;
  wire L111P_0a;
  wire [31:0] L111A_0r0;
  wire [31:0] L111A_0r1;
  wire L111A_0a;
  wire L112P_0r;
  wire L112P_0a;
  wire L112A_0r;
  wire L112A_0a;
  wire [31:0] L113_0r0;
  wire [31:0] L113_0r1;
  wire L113_0a;
  wire [63:0] L114P_0r0;
  wire [63:0] L114P_0r1;
  wire L114P_0a;
  wire [63:0] L114A_0r0;
  wire [63:0] L114A_0r1;
  wire L114A_0a;
  wire [32:0] L115_0r0;
  wire [32:0] L115_0r1;
  wire L115_0a;
  wire L116P_0r;
  wire L116P_0a;
  wire L116A_0r;
  wire L116A_0a;
  wire L120P_0r;
  wire L120P_0a;
  wire L120A_0r;
  wire L120A_0a;
  wire [32:0] L125P_0r0;
  wire [32:0] L125P_0r1;
  wire L125P_0a;
  wire [32:0] L125A_0r0;
  wire [32:0] L125A_0r1;
  wire L125A_0a;
  wire L128P_0r;
  wire L128P_0a;
  wire L128A_0r;
  wire L128A_0a;
  wire L131P_0r;
  wire L131P_0a;
  wire L131A_0r;
  wire L131A_0a;
  wire L136_0r0;
  wire L136_0r1;
  wire L136_0a;
  wire L138_0r;
  wire L138_0a;
  wire L140_0r;
  wire L140_0a;
  wire L143_0r;
  wire L143_0a;
  wire L145P_0r;
  wire L145P_0a;
  wire L145A_0r;
  wire L145A_0a;
  wire L148P_0r;
  wire L148P_0a;
  wire L148A_0r;
  wire L148A_0a;
  wire [2:0] L149P_0r0;
  wire [2:0] L149P_0r1;
  wire L149P_0a;
  wire [2:0] L149A_0r0;
  wire [2:0] L149A_0r1;
  wire L149A_0a;
  wire L150P_0r;
  wire L150P_0a;
  wire L150A_0r;
  wire L150A_0a;
  wire L151P_0r;
  wire L151P_0a;
  wire L151A_0r;
  wire L151A_0a;
  wire [2:0] L152P_0r0;
  wire [2:0] L152P_0r1;
  wire L152P_0a;
  wire [2:0] L152A_0r0;
  wire [2:0] L152A_0r1;
  wire L152A_0a;
  wire L153P_0r;
  wire L153P_0a;
  wire L153A_0r;
  wire L153A_0a;
  wire [2:0] L154P_0r0;
  wire [2:0] L154P_0r1;
  wire L154P_0a;
  wire [2:0] L154A_0r0;
  wire [2:0] L154A_0r1;
  wire L154A_0a;
  wire L155_0r;
  wire L155_0a;
  wire [2:0] L156P_0r0;
  wire [2:0] L156P_0r1;
  wire L156P_0a;
  wire [2:0] L156A_0r0;
  wire [2:0] L156A_0r1;
  wire L156A_0a;
  wire [2:0] L157P_0r0;
  wire [2:0] L157P_0r1;
  wire L157P_0a;
  wire [2:0] L157A_0r0;
  wire [2:0] L157A_0r1;
  wire L157A_0a;
  wire [2:0] L158P_0r0;
  wire [2:0] L158P_0r1;
  wire L158P_0a;
  wire [2:0] L158A_0r0;
  wire [2:0] L158A_0r1;
  wire L158A_0a;
  wire [2:0] L159_0r0;
  wire [2:0] L159_0r1;
  wire L159_0a;
  wire [2:0] L160P_0r0;
  wire [2:0] L160P_0r1;
  wire L160P_0a;
  wire [2:0] L160A_0r0;
  wire [2:0] L160A_0r1;
  wire L160A_0a;
  wire [2:0] L161P_0r0;
  wire [2:0] L161P_0r1;
  wire L161P_0a;
  wire [2:0] L161A_0r0;
  wire [2:0] L161A_0r1;
  wire L161A_0a;
  wire [31:0] L162P_0r0;
  wire [31:0] L162P_0r1;
  wire L162P_0a;
  wire [31:0] L162A_0r0;
  wire [31:0] L162A_0r1;
  wire L162A_0a;
  wire L163P_0r;
  wire L163P_0a;
  wire L163A_0r;
  wire L163A_0a;
  wire L164_0r;
  wire L164_0a;
  wire [31:0] L165P_0r0;
  wire [31:0] L165P_0r1;
  wire L165P_0a;
  wire [31:0] L165A_0r0;
  wire [31:0] L165A_0r1;
  wire L165A_0a;
  wire L166_0r;
  wire L166_0a;
  wire [31:0] L167P_0r0;
  wire [31:0] L167P_0r1;
  wire L167P_0a;
  wire [31:0] L167A_0r0;
  wire [31:0] L167A_0r1;
  wire L167A_0a;
  wire L168_0r;
  wire L168_0a;
  wire [31:0] L169_0r0;
  wire [31:0] L169_0r1;
  wire L169_0a;
  wire [2:0] L170P_0r0;
  wire [2:0] L170P_0r1;
  wire L170P_0a;
  wire [2:0] L170A_0r0;
  wire [2:0] L170A_0r1;
  wire L170A_0a;
  wire [2:0] L171P_0r0;
  wire [2:0] L171P_0r1;
  wire L171P_0a;
  wire [2:0] L171A_0r0;
  wire [2:0] L171A_0r1;
  wire L171A_0a;
  wire [2:0] L172P_0r0;
  wire [2:0] L172P_0r1;
  wire L172P_0a;
  wire [2:0] L172A_0r0;
  wire [2:0] L172A_0r1;
  wire L172A_0a;
  wire [2:0] L173P_0r0;
  wire [2:0] L173P_0r1;
  wire L173P_0a;
  wire [2:0] L173A_0r0;
  wire [2:0] L173A_0r1;
  wire L173A_0a;
  wire [2:0] L174P_0r0;
  wire [2:0] L174P_0r1;
  wire L174P_0a;
  wire [2:0] L174A_0r0;
  wire [2:0] L174A_0r1;
  wire L174A_0a;
  wire [31:0] L175P_0r0;
  wire [31:0] L175P_0r1;
  wire L175P_0a;
  wire [31:0] L175A_0r0;
  wire [31:0] L175A_0r1;
  wire L175A_0a;
  wire L176P_0r;
  wire L176P_0a;
  wire L176A_0r;
  wire L176A_0a;
  wire L177P_0r;
  wire L177P_0a;
  wire L177A_0r;
  wire L177A_0a;
  wire [31:0] L178P_0r0;
  wire [31:0] L178P_0r1;
  wire L178P_0a;
  wire [31:0] L178A_0r0;
  wire [31:0] L178A_0r1;
  wire L178A_0a;
  wire L179_0r;
  wire L179_0a;
  wire [31:0] L180P_0r0;
  wire [31:0] L180P_0r1;
  wire L180P_0a;
  wire [31:0] L180A_0r0;
  wire [31:0] L180A_0r1;
  wire L180A_0a;
  wire [1:0] L181P_0r0;
  wire [1:0] L181P_0r1;
  wire L181P_0a;
  wire [1:0] L181A_0r0;
  wire [1:0] L181A_0r1;
  wire L181A_0a;
  wire [1:0] L182_0r0;
  wire [1:0] L182_0r1;
  wire L182_0a;
  wire [1:0] L183P_0r0;
  wire [1:0] L183P_0r1;
  wire L183P_0a;
  wire [1:0] L183A_0r0;
  wire [1:0] L183A_0r1;
  wire L183A_0a;
  wire [1:0] L184P_0r0;
  wire [1:0] L184P_0r1;
  wire L184P_0a;
  wire [1:0] L184A_0r0;
  wire [1:0] L184A_0r1;
  wire L184A_0a;
  wire [31:0] L185P_0r0;
  wire [31:0] L185P_0r1;
  wire L185P_0a;
  wire [31:0] L185A_0r0;
  wire [31:0] L185A_0r1;
  wire L185A_0a;
  wire L186P_0r;
  wire L186P_0a;
  wire L186A_0r;
  wire L186A_0a;
  wire L187P_0r;
  wire L187P_0a;
  wire L187A_0r;
  wire L187A_0a;
  wire [31:0] L188P_0r0;
  wire [31:0] L188P_0r1;
  wire L188P_0a;
  wire [31:0] L188A_0r0;
  wire [31:0] L188A_0r1;
  wire L188A_0a;
  wire L189P_0r;
  wire L189P_0a;
  wire L189A_0r;
  wire L189A_0a;
  wire [31:0] L190_0r0;
  wire [31:0] L190_0r1;
  wire L190_0a;
  wire L191_0r;
  wire L191_0a;
  wire [31:0] L192_0r0;
  wire [31:0] L192_0r1;
  wire L192_0a;
  wire [2:0] L193P_0r0;
  wire [2:0] L193P_0r1;
  wire L193P_0a;
  wire [2:0] L193A_0r0;
  wire [2:0] L193A_0r1;
  wire L193A_0a;
  wire [2:0] L194P_0r0;
  wire [2:0] L194P_0r1;
  wire L194P_0a;
  wire [2:0] L194A_0r0;
  wire [2:0] L194A_0r1;
  wire L194A_0a;
  wire [2:0] L195_0r0;
  wire [2:0] L195_0r1;
  wire L195_0a;
  wire [2:0] L196P_0r0;
  wire [2:0] L196P_0r1;
  wire L196P_0a;
  wire [2:0] L196A_0r0;
  wire [2:0] L196A_0r1;
  wire L196A_0a;
  wire [2:0] L197P_0r0;
  wire [2:0] L197P_0r1;
  wire L197P_0a;
  wire [2:0] L197A_0r0;
  wire [2:0] L197A_0r1;
  wire L197A_0a;
  wire L198P_0r;
  wire L198P_0a;
  wire L198A_0r;
  wire L198A_0a;
  wire [31:0] L199_0r0;
  wire [31:0] L199_0r1;
  wire L199_0a;
  wire L200_0r;
  wire L200_0a;
  wire [63:0] L206_0r0;
  wire [63:0] L206_0r1;
  wire L206_0a;
  wire [31:0] L211_0r0;
  wire [31:0] L211_0r1;
  wire L211_0a;
  wire L216_0r;
  wire L216_0a;
  wire L217_0r;
  wire L217_0a;
  wire L218_0r;
  wire L218_0a;
  wire [63:0] L224_0r0;
  wire [63:0] L224_0r1;
  wire L224_0a;
  wire [31:0] L229_0r0;
  wire [31:0] L229_0r1;
  wire L229_0a;
  wire L234_0r;
  wire L234_0a;
  wire L235_0r;
  wire L235_0a;
  wire L236_0r;
  wire L236_0a;
  wire [63:0] L242_0r0;
  wire [63:0] L242_0r1;
  wire L242_0a;
  wire [31:0] L247_0r0;
  wire [31:0] L247_0r1;
  wire L247_0a;
  wire [31:0] L249_0r0;
  wire [31:0] L249_0r1;
  wire L249_0a;
  wire L252_0r;
  wire L252_0a;
  wire L253P_0r;
  wire L253P_0a;
  wire L253A_0r;
  wire L253A_0a;
  wire L254_0r;
  wire L254_0a;
  wire L255P_0r;
  wire L255P_0a;
  wire L255A_0r;
  wire L255A_0a;
  wire L257P_0r;
  wire L257P_0a;
  wire L257A_0r;
  wire L257A_0a;
  wire L260P_0r;
  wire L260P_0a;
  wire L260A_0r;
  wire L260A_0a;
  wire [31:0] L264P_0r0;
  wire [31:0] L264P_0r1;
  wire L264P_0a;
  wire [31:0] L264A_0r0;
  wire [31:0] L264A_0r1;
  wire L264A_0a;
  wire L267_0r;
  wire L267_0a;
  wire [32:0] L272P_0r0;
  wire [32:0] L272P_0r1;
  wire L272P_0a;
  wire [32:0] L272A_0r0;
  wire [32:0] L272A_0r1;
  wire L272A_0a;
  wire L275P_0r;
  wire L275P_0a;
  wire L275A_0r;
  wire L275A_0a;
  wire L277P_0r;
  wire L277P_0a;
  wire L277A_0r;
  wire L277A_0a;
  wire L278_0r;
  wire L278_0a;
  wire L281P_0r;
  wire L281P_0a;
  wire L281A_0r;
  wire L281A_0a;
  wire L284P_0r;
  wire L284P_0a;
  wire L284A_0r;
  wire L284A_0a;
  wire [31:0] L286_0r0;
  wire [31:0] L286_0r1;
  wire L286_0a;
  wire [31:0] L288_0r0;
  wire [31:0] L288_0r1;
  wire L288_0a;
  wire [2:0] L289_0r0;
  wire [2:0] L289_0r1;
  wire L289_0a;
  wire [2:0] L290_0r0;
  wire [2:0] L290_0r1;
  wire L290_0a;
  wire [2:0] L291_0r0;
  wire [2:0] L291_0r1;
  wire L291_0a;
  wire [2:0] L292_0r0;
  wire [2:0] L292_0r1;
  wire L292_0a;
  wire [34:0] L293_0r0;
  wire [34:0] L293_0r1;
  wire L293_0a;
  wire [31:0] L295_0r0;
  wire [31:0] L295_0r1;
  wire L295_0a;
  wire [31:0] L297_0r0;
  wire [31:0] L297_0r1;
  wire L297_0a;
  wire [31:0] L299_0r0;
  wire [31:0] L299_0r1;
  wire L299_0a;
  wire [31:0] L302P_0r0;
  wire [31:0] L302P_0r1;
  wire L302P_0a;
  wire [31:0] L302A_0r0;
  wire [31:0] L302A_0r1;
  wire L302A_0a;
  wire [31:0] L308P_0r0;
  wire [31:0] L308P_0r1;
  wire L308P_0a;
  wire [31:0] L308A_0r0;
  wire [31:0] L308A_0r1;
  wire L308A_0a;
  wire L309_0r;
  wire L309_0a;
  wire L310_0r;
  wire L310_0a;
  wire [31:0] L311_0r0;
  wire [31:0] L311_0r1;
  wire L311_0a;
  wire L312_0r;
  wire L312_0a;
  wire [31:0] L313P_0r0;
  wire [31:0] L313P_0r1;
  wire L313P_0a;
  wire [31:0] L313A_0r0;
  wire [31:0] L313A_0r1;
  wire L313A_0a;
  wire [1:0] L314_0r0;
  wire [1:0] L314_0r1;
  wire L314_0a;
  wire [1:0] L315_0r0;
  wire [1:0] L315_0r1;
  wire L315_0a;
  wire [1:0] L316_0r0;
  wire [1:0] L316_0r1;
  wire L316_0a;
  wire [1:0] L317P_0r0;
  wire [1:0] L317P_0r1;
  wire L317P_0a;
  wire [1:0] L317A_0r0;
  wire [1:0] L317A_0r1;
  wire L317A_0a;
  wire [31:0] L318P_0r0;
  wire [31:0] L318P_0r1;
  wire L318P_0a;
  wire [31:0] L318A_0r0;
  wire [31:0] L318A_0r1;
  wire L318A_0a;
  wire L319P_0r;
  wire L319P_0a;
  wire L319A_0r;
  wire L319A_0a;
  wire L320P_0r;
  wire L320P_0a;
  wire L320A_0r;
  wire L320A_0a;
  wire [31:0] L321_0r0;
  wire [31:0] L321_0r1;
  wire L321_0a;
  wire L322_0r;
  wire L322_0a;
  wire [31:0] L323_0r0;
  wire [31:0] L323_0r1;
  wire L323_0a;
  wire [1:0] L324P_0r0;
  wire [1:0] L324P_0r1;
  wire L324P_0a;
  wire [1:0] L324A_0r0;
  wire [1:0] L324A_0r1;
  wire L324A_0a;
  wire [1:0] L325_0r0;
  wire [1:0] L325_0r1;
  wire L325_0a;
  wire [1:0] L326P_0r0;
  wire [1:0] L326P_0r1;
  wire L326P_0a;
  wire [1:0] L326A_0r0;
  wire [1:0] L326A_0r1;
  wire L326A_0a;
  wire [1:0] L327P_0r0;
  wire [1:0] L327P_0r1;
  wire L327P_0a;
  wire [1:0] L327A_0r0;
  wire [1:0] L327A_0r1;
  wire L327A_0a;
  wire [1:0] L332_0r0;
  wire [1:0] L332_0r1;
  wire L332_0a;
  wire [1:0] L333P_0r0;
  wire [1:0] L333P_0r1;
  wire L333P_0a;
  wire [1:0] L333A_0r0;
  wire [1:0] L333A_0r1;
  wire L333A_0a;
  wire [1:0] L334P_0r0;
  wire [1:0] L334P_0r1;
  wire L334P_0a;
  wire [1:0] L334A_0r0;
  wire [1:0] L334A_0r1;
  wire L334A_0a;
  wire [33:0] L335_0r0;
  wire [33:0] L335_0r1;
  wire L335_0a;
  wire L338P_0r;
  wire L338P_0a;
  wire L338A_0r;
  wire L338A_0a;
  wire L345P_0r0;
  wire L345P_0r1;
  wire L345P_0a;
  wire L345A_0r0;
  wire L345A_0r1;
  wire L345A_0a;
  wire L346P_0r0;
  wire L346P_0r1;
  wire L346P_0a;
  wire L346A_0r0;
  wire L346A_0r1;
  wire L346A_0a;
  wire [2:0] L347P_0r0;
  wire [2:0] L347P_0r1;
  wire L347P_0a;
  wire [2:0] L347A_0r0;
  wire [2:0] L347A_0r1;
  wire L347A_0a;
  wire L348P_0r0;
  wire L348P_0r1;
  wire L348P_0a;
  wire L348A_0r0;
  wire L348A_0r1;
  wire L348A_0a;
  wire [2:0] L349_0r0;
  wire [2:0] L349_0r1;
  wire L349_0a;
  wire [31:0] L350_0r0;
  wire [31:0] L350_0r1;
  wire L350_0a;
  wire [31:0] L351_0r0;
  wire [31:0] L351_0r1;
  wire L351_0a;
  wire [2:0] L352_0r0;
  wire [2:0] L352_0r1;
  wire L352_0a;
  wire [31:0] L353P_0r0;
  wire [31:0] L353P_0r1;
  wire L353P_0a;
  wire [31:0] L353A_0r0;
  wire [31:0] L353A_0r1;
  wire L353A_0a;
  wire L355_0r;
  wire L355_0a;
  wire L356_0r;
  wire L356_0a;
  wire L357_0r;
  wire L357_0a;
  wire [31:0] L358P_0r0;
  wire [31:0] L358P_0r1;
  wire L358P_0a;
  wire [31:0] L358A_0r0;
  wire [31:0] L358A_0r1;
  wire L358A_0a;
  wire [31:0] L359P_0r0;
  wire [31:0] L359P_0r1;
  wire L359P_0a;
  wire [31:0] L359A_0r0;
  wire [31:0] L359A_0r1;
  wire L359A_0a;
  wire [31:0] L360P_0r0;
  wire [31:0] L360P_0r1;
  wire L360P_0a;
  wire [31:0] L360A_0r0;
  wire [31:0] L360A_0r1;
  wire L360A_0a;
  wire L361P_0r;
  wire L361P_0a;
  wire L361A_0r;
  wire L361A_0a;
  wire L362P_0r;
  wire L362P_0a;
  wire L362A_0r;
  wire L362A_0a;
  wire L363P_0r;
  wire L363P_0a;
  wire L363A_0r;
  wire L363A_0a;
  wire L364P_0r;
  wire L364P_0a;
  wire L364A_0r;
  wire L364A_0a;
  wire L366P_0r;
  wire L366P_0a;
  wire L366A_0r;
  wire L366A_0a;
  wire L367P_0r;
  wire L367P_0a;
  wire L367A_0r;
  wire L367A_0a;
  wire L385P_0r;
  wire L385P_0a;
  wire L385A_0r;
  wire L385A_0a;
  wire [31:0] L395P_0r0;
  wire [31:0] L395P_0r1;
  wire L395P_0a;
  wire [31:0] L395A_0r0;
  wire [31:0] L395A_0r1;
  wire L395A_0a;
  tko0m32_1nm32b1 I0 (L355_0r, L355_0a, L313A_0r0[31:0], L313A_0r1[31:0], L313A_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I1 (L14P_0r, L14P_0a, L7_0r, L7_0a, L312_0r, L312_0a, L355_0r, L355_0a, reset);
  tkj0m0_0 I2 (L9_0r, L9_0a, L13P_0r, L13P_0a, L277A_0r, L277A_0a, reset);
  tko0m32_1nm32b0 I3 (L356_0r, L356_0a, L192_0r0[31:0], L192_0r1[31:0], L192_0a, reset);
  tko0m3_1nm3b0 I4 (L357_0r, L357_0a, L156A_0r0[2:0], L156A_0r1[2:0], L156A_0a, reset);
  tko32m32_1nm32b0_2subt1o0w32bi0w32b I5 (L358P_0r0[31:0], L358P_0r1[31:0], L358P_0a, L178A_0r0[31:0], L178A_0r1[31:0], L178A_0a, reset);
  tkf4mo0w0_o0w3 I6 (L68_0r0[3:0], L68_0r1[3:0], L68_0a, L153A_0r, L153A_0a, L154A_0r0[2:0], L154A_0r1[2:0], L154A_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I7 (L72P_0r, L72P_0a, L63A_0r, L63A_0a, L362A_0r, L362A_0a, L177A_0r, L177A_0a, reset);
  tkj0m0_0 I8 (L61_0r, L61_0a, L71_0r, L71_0a, L73A_0r, L73A_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I9 (L54_0r0, L54_0r1, L54_0a, L56A_0r, L56A_0a, L72A_0r, L72A_0a, reset);
  tkm2x0b I10 (L56P_0r, L56P_0a, L73P_0r, L73P_0a, L75A_0r, L75A_0a, reset);
  tko32m32_1nm32b0_2subt1o0w32bi0w32b I11 (L359P_0r0[31:0], L359P_0r1[31:0], L359P_0a, L167A_0r0[31:0], L167A_0r1[31:0], L167A_0a, reset);
  tkf4mo0w0_o0w3 I12 (L94P_0r0[3:0], L94P_0r1[3:0], L94P_0a, L151A_0r, L151A_0a, L152A_0r0[2:0], L152A_0r1[2:0], L152A_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I13 (L98P_0r, L98P_0a, L89A_0r, L89A_0a, L361A_0r, L361A_0a, L166_0r, L166_0a, reset);
  tkj0m0_0 I14 (L87_0r, L87_0a, L97_0r, L97_0a, L99A_0r, L99A_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I15 (L80_0r0, L80_0r1, L80_0a, L82A_0r, L82A_0a, L98A_0r, L98A_0a, reset);
  tkj64m32_32 I16 (L111P_0r0[31:0], L111P_0r1[31:0], L111P_0a, L113_0r0[31:0], L113_0r1[31:0], L113_0a, L114A_0r0[63:0], L114A_0r1[63:0], L114A_0a, reset);
  tko64m33_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b I17 (L114P_0r0[63:0], L114P_0r1[63:0], L114P_0a, L115_0r0[32:0], L115_0r1[32:0], L115_0a, reset);
  tkf33mo0w0_o0w32 I18 (L115_0r0[32:0], L115_0r1[32:0], L115_0a, L189A_0r, L189A_0a, L190_0r0[31:0], L190_0r1[31:0], L190_0a, reset);
  tkf0mo0w0_o0w0 I19 (L116P_0r, L116P_0a, L110A_0r, L110A_0a, L112A_0r, L112A_0a, reset);
  tkf33mo0w0_o0w32 I20 (L125P_0r0[32:0], L125P_0r1[32:0], L125P_0a, L164_0r, L164_0a, L165A_0r0[31:0], L165A_0r1[31:0], L165A_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I21 (L106_0r0, L106_0r1, L106_0a, L131A_0r, L131A_0a, L116A_0r, L116A_0a, reset);
  tkm3x0b I22 (L82P_0r, L82P_0a, L99P_0r, L99P_0a, L128P_0r, L128P_0a, L101A_0r, L101A_0a, reset);
  tko32m32_1nm32b0_2subt1o0w32bi0w32b I23 (L360P_0r0[31:0], L360P_0r1[31:0], L360P_0a, L188A_0r0[31:0], L188A_0r1[31:0], L188A_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I24 (L136_0r0, L136_0r1, L136_0a, L138_0r, L138_0a, L140_0r, L140_0a, reset);
  tkm2x0b I25 (L138_0r, L138_0a, L143_0r, L143_0a, L145A_0r, L145A_0a, reset);
  tkf0mo0w0_o0w0 I26 (L45_0r, L45_0a, L155_0r, L155_0a, L357_0r, L357_0a, reset);
  tkm3x3b I27 (L152P_0r0[2:0], L152P_0r1[2:0], L152P_0a, L154P_0r0[2:0], L154P_0r1[2:0], L154P_0a, L156P_0r0[2:0], L156P_0r1[2:0], L156P_0a, L149A_0r0[2:0], L149A_0r1[2:0], L149A_0a, reset);
  tko0m3_1nm3b1 I28 (L151P_0r, L151P_0a, L157A_0r0[2:0], L157A_0r1[2:0], L157A_0a, reset);
  tko0m3_1nm3b2 I29 (L153P_0r, L153P_0a, L158A_0r0[2:0], L158A_0r1[2:0], L158A_0a, reset);
  tko0m3_1nm3b4 I30 (L155_0r, L155_0a, L159_0r0[2:0], L159_0r1[2:0], L159_0a, reset);
  tkm3x3b I31 (L157P_0r0[2:0], L157P_0r1[2:0], L157P_0a, L158P_0r0[2:0], L158P_0r1[2:0], L158P_0a, L159_0r0[2:0], L159_0r1[2:0], L159_0a, L160A_0r0[2:0], L160A_0r1[2:0], L160A_0a, reset);
  tkj3m0_3 I32 (L150P_0r, L150P_0a, L160P_0r0[2:0], L160P_0r1[2:0], L160P_0a, L161A_0r0[2:0], L161A_0r1[2:0], L161A_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I33 (L161P_0r0[2:0], L161P_0r1[2:0], L161P_0a, L97_0r, L97_0a, L71_0r, L71_0a, L49A_0r, L49A_0a, reset);
  tkvneg3_wo0w3_ro0w3o0w3o0w3 I34 (L149P_0r0[2:0], L149P_0r1[2:0], L149P_0a, L150A_0r, L150A_0a, L131P_0r, L131P_0a, L89P_0r, L89P_0a, L63P_0r, L63P_0a, L352_0r0[2:0], L352_0r1[2:0], L352_0a, L349_0r0[2:0], L349_0r1[2:0], L349_0a, L347A_0r0[2:0], L347A_0r1[2:0], L347A_0a, reset);
  tkm3x32b I35 (L165P_0r0[31:0], L165P_0r1[31:0], L165P_0a, L167P_0r0[31:0], L167P_0r1[31:0], L167P_0a, L169_0r0[31:0], L169_0r1[31:0], L169_0a, L162A_0r0[31:0], L162A_0r1[31:0], L162A_0a, reset);
  tko0m3_1nm3b1 I36 (L164_0r, L164_0a, L170A_0r0[2:0], L170A_0r1[2:0], L170A_0a, reset);
  tko0m3_1nm3b2 I37 (L166_0r, L166_0a, L171A_0r0[2:0], L171A_0r1[2:0], L171A_0a, reset);
  tko0m3_1nm3b4 I38 (L168_0r, L168_0a, L172A_0r0[2:0], L172A_0r1[2:0], L172A_0a, reset);
  tkm3x3b I39 (L170P_0r0[2:0], L170P_0r1[2:0], L170P_0a, L171P_0r0[2:0], L171P_0r1[2:0], L171P_0a, L172P_0r0[2:0], L172P_0r1[2:0], L172P_0a, L173A_0r0[2:0], L173A_0r1[2:0], L173A_0a, reset);
  tkj3m0_3 I40 (L163P_0r, L163P_0a, L173P_0r0[2:0], L173P_0r1[2:0], L173P_0a, L174A_0r0[2:0], L174A_0r1[2:0], L174A_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I41 (L174P_0r0[2:0], L174P_0r1[2:0], L174P_0a, L128A_0r, L128A_0a, L87_0r, L87_0a, L38_0r, L38_0a, reset);
  tkvr332_wo0w32_ro0w32o0w32o0w32o31w1 I42 (L162P_0r0[31:0], L162P_0r1[31:0], L162P_0a, L163A_0r, L163A_0a, L120P_0r, L120P_0a, L101P_0r, L101P_0a, L361P_0r, L361P_0a, L75P_0r, L75P_0a, L351_0r0[31:0], L351_0r1[31:0], L351_0a, L350_0r0[31:0], L350_0r1[31:0], L350_0a, L359A_0r0[31:0], L359A_0r1[31:0], L359A_0a, L348A_0r0, L348A_0r1, L348A_0a, reset);
  tkf32mo0w0_o0w32 I43 (L39_0r0[31:0], L39_0r1[31:0], L39_0a, L179_0r, L179_0a, L180A_0r0[31:0], L180A_0r1[31:0], L180A_0a, reset);
  tkm2x32b I44 (L178P_0r0[31:0], L178P_0r1[31:0], L178P_0a, L180P_0r0[31:0], L180P_0r1[31:0], L180P_0a, L175A_0r0[31:0], L175A_0r1[31:0], L175A_0a, reset);
  tko0m2_1nm2b1 I45 (L177P_0r, L177P_0a, L181A_0r0[1:0], L181A_0r1[1:0], L181A_0a, reset);
  tko0m2_1nm2b2 I46 (L179_0r, L179_0a, L182_0r0[1:0], L182_0r1[1:0], L182_0a, reset);
  tkm2x2b I47 (L181P_0r0[1:0], L181P_0r1[1:0], L181P_0a, L182_0r0[1:0], L182_0r1[1:0], L182_0a, L183A_0r0[1:0], L183A_0r1[1:0], L183A_0a, reset);
  tkj2m0_2 I48 (L176P_0r, L176P_0a, L183P_0r0[1:0], L183P_0r1[1:0], L183P_0a, L184A_0r0[1:0], L184A_0r1[1:0], L184A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I49 (L184P_0r0[1:0], L184P_0r1[1:0], L184P_0a, L61_0r, L61_0a, L41_0r, L41_0a, reset);
  tkvr232_wo0w32_ro0w32o0w32o31w1 I50 (L175P_0r0[31:0], L175P_0r1[31:0], L175P_0a, L176A_0r, L176A_0a, L112P_0r, L112P_0a, L362P_0r, L362P_0a, L49P_0r, L49P_0a, L113_0r0[31:0], L113_0r1[31:0], L113_0a, L358A_0r0[31:0], L358A_0r1[31:0], L358A_0a, L346A_0r0, L346A_0r1, L346A_0a, reset);
  tkf0mo0w0_o0w0 I51 (L41_0r, L41_0a, L191_0r, L191_0a, L356_0r, L356_0a, reset);
  tkm3x32b I52 (L188P_0r0[31:0], L188P_0r1[31:0], L188P_0a, L190_0r0[31:0], L190_0r1[31:0], L190_0a, L192_0r0[31:0], L192_0r1[31:0], L192_0a, L185A_0r0[31:0], L185A_0r1[31:0], L185A_0a, reset);
  tko0m3_1nm3b1 I53 (L187P_0r, L187P_0a, L193A_0r0[2:0], L193A_0r1[2:0], L193A_0a, reset);
  tko0m3_1nm3b2 I54 (L189P_0r, L189P_0a, L194A_0r0[2:0], L194A_0r1[2:0], L194A_0a, reset);
  tko0m3_1nm3b4 I55 (L191_0r, L191_0a, L195_0r0[2:0], L195_0r1[2:0], L195_0a, reset);
  tkm3x3b I56 (L193P_0r0[2:0], L193P_0r1[2:0], L193P_0a, L194P_0r0[2:0], L194P_0r1[2:0], L194P_0a, L195_0r0[2:0], L195_0r1[2:0], L195_0a, L196A_0r0[2:0], L196A_0r1[2:0], L196A_0a, reset);
  tkj3m0_3 I57 (L186P_0r, L186P_0a, L196P_0r0[2:0], L196P_0r1[2:0], L196P_0a, L197A_0r0[2:0], L197A_0r1[2:0], L197A_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I58 (L197P_0r0[2:0], L197P_0r1[2:0], L197P_0a, L143_0r, L143_0a, L120A_0r, L120A_0a, L45_0r, L45_0a, reset);
  tkvr132_wo0w32_ro0w32o0w32o0w32 I59 (L185P_0r0[31:0], L185P_0r1[31:0], L185P_0a, L186A_0r, L186A_0a, L366P_0r, L366P_0a, L363P_0r, L363P_0a, L110P_0r, L110P_0a, L288_0r0[31:0], L288_0r1[31:0], L288_0a, L360A_0r0[31:0], L360A_0r1[31:0], L360A_0a, L111A_0r0[31:0], L111A_0r1[31:0], L111A_0a, reset);
  tkf0mo0w0_o0w0 I60 (L218_0r, L218_0a, L216_0r, L216_0a, L217_0r, L217_0a, reset);
  tkf0mo0w0_o0w0 I61 (L236_0r, L236_0a, L234_0r, L234_0a, L235_0r, L235_0a, reset);
  tkf0mo0w0_o0w0 I62 (L254_0r, L254_0a, L252_0r, L252_0a, L253A_0r, L253A_0a, reset);
  tks32_o0w32_3cfffffffcm4cfffffff8m5cfffffff8m6cfffffff8m8cfffffff0m9cfffffff0macfffffff0m10cffffffe0m11cffffffe0m12cffffffe0m20cffffffc0m21cffffffc0m22cffffffc0m40cffffff80m41cffffff80m42cffffff80m80cffffff00m81cffffff00m82cffffff00m100cfffffe00m101cfffffe00m102cfffffe00m200cfffffc00m201cfffffc00m202cfffffc00m400cfffff800m401cfffff800m402cfffff800m800cfffff000m801cfffff000m802cfffff000m1000cffffe000m1001cffffe000m1002cffffe000m2000cffffc000m2001cffffc000m2002cffffc000m4000cffff8000m4001cffff8000m4002cffff8000m8000cffff0000m8001cffff0000m8002cffff0000m10000cfffe0000m10001cfffe0000m10002cfffe0000m20000cfffc0000m20001cfffc0000m20002cfffc0000m40000cfff80000m40001cfff80000m40002cfff80000m80000cfff00000m80001cfff00000m80002cfff00000m100000cffe00000m100001cffe00000m100002cffe00000m200000cffc00000m200001cffc00000m200002cffc00000m400000cff800000m400001cff800000m400002cff800000m800000cff000000m800001cff000000m800002cff000000m1000000cfe000000m1000001cfe000000m1000002cfe000000m2000000cfc000000m2000001cfc000000m2000002cfc000000m4000000cf8000000m4000001cf8000000m4000002cf8000000m8000000cf0000000m8000001cf0000000m8000002cf0000000m10000000ce0000000m10000001ce0000000m10000002ce0000000m20000000cc0000000m20000001cc0000000m20000002cc0000000m40000000c80000000m40000001c80000000m40000002c80000000m80000000m80000001m80000002o0w0_0o0w0_1o0w0_2o0w0 I63 (L199_0r0[31:0], L199_0r1[31:0], L199_0a, L200_0r, L200_0a, L218_0r, L218_0a, L236_0r, L236_0a, L254_0r, L254_0a, reset);
  tkm2x0b I64 (L338P_0r, L338P_0a, L200_0r, L200_0a, L255A_0r, L255A_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0 I65 (L260P_0r, L260P_0a, L257A_0r, L257A_0a, L385A_0r, L385A_0a, L168_0r, L168_0a, L364A_0r, L364A_0a, L198A_0r, L198A_0a, reset);
  tkf33mo0w0_o0w32 I66 (L272P_0r0[32:0], L272P_0r1[32:0], L272P_0a, L310_0r, L310_0a, L311_0r0[31:0], L311_0r1[31:0], L311_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I67 (L21_0r0, L21_0r1, L21_0a, L278_0r, L278_0a, L260A_0r, L260A_0a, reset);
  tkm2x0b I68 (L277P_0r, L277P_0a, L275P_0r, L275P_0a, L16A_0r, L16A_0a, reset);
  tkj32m32_0 I69 (L286_0r0[31:0], L286_0r1[31:0], L286_0a, L38_0r, L38_0a, L39_0r0[31:0], L39_0r1[31:0], L39_0a, reset);
  tko0m3_1nm3b1 I70 (L216_0r, L216_0a, L289_0r0[2:0], L289_0r1[2:0], L289_0a, reset);
  tko0m3_1nm3b2 I71 (L234_0r, L234_0a, L290_0r0[2:0], L290_0r1[2:0], L290_0a, reset);
  tko0m3_1nm3b4 I72 (L252_0r, L252_0a, L291_0r0[2:0], L291_0r1[2:0], L291_0a, reset);
  tkm3x3b I73 (L289_0r0[2:0], L289_0r1[2:0], L289_0a, L290_0r0[2:0], L290_0r1[2:0], L290_0a, L291_0r0[2:0], L291_0r1[2:0], L291_0a, L292_0r0[2:0], L292_0r1[2:0], L292_0a, reset);
  tkj35m32_3 I74 (L288_0r0[31:0], L288_0r1[31:0], L288_0a, L292_0r0[2:0], L292_0r1[2:0], L292_0a, L293_0r0[34:0], L293_0r1[34:0], L293_0a, reset);
  tks35_o32w3_1o0w32_2o0w32_4o0w32 I75 (L293_0r0[34:0], L293_0r1[34:0], L293_0a, L211_0r0[31:0], L211_0r1[31:0], L211_0a, L229_0r0[31:0], L229_0r1[31:0], L229_0a, L247_0r0[31:0], L247_0r1[31:0], L247_0a, reset);
  tkvxV32_wo0w32_ro0w32 I76 (L4P_0r0[31:0], L4P_0r1[31:0], L4P_0a, L14A_0r, L14A_0a, L364P_0r, L364P_0a, L286_0r0[31:0], L286_0r1[31:0], L286_0a, reset);
  tkm2x32b I77 (L311_0r0[31:0], L311_0r1[31:0], L311_0a, L313P_0r0[31:0], L313P_0r1[31:0], L313P_0a, L308A_0r0[31:0], L308A_0r1[31:0], L308A_0a, reset);
  tko0m2_1nm2b1 I78 (L310_0r, L310_0a, L314_0r0[1:0], L314_0r1[1:0], L314_0a, reset);
  tko0m2_1nm2b2 I79 (L312_0r, L312_0a, L315_0r0[1:0], L315_0r1[1:0], L315_0a, reset);
  tkm2x2b I80 (L314_0r0[1:0], L314_0r1[1:0], L314_0a, L315_0r0[1:0], L315_0r1[1:0], L315_0a, L316_0r0[1:0], L316_0r1[1:0], L316_0a, reset);
  tkj2m0_2 I81 (L309_0r, L309_0a, L316_0r0[1:0], L316_0r1[1:0], L316_0a, L317A_0r0[1:0], L317A_0r1[1:0], L317A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I82 (L317P_0r0[1:0], L317P_0r1[1:0], L317P_0a, L275A_0r, L275A_0a, L13A_0r, L13A_0a, reset);
  tkvi32_wo0w32_ro0w32o0w32o31w1 I83 (L308P_0r0[31:0], L308P_0r1[31:0], L308P_0a, L309_0r, L309_0a, L267_0r, L267_0a, L198P_0r, L198P_0a, L16P_0r, L16P_0a, L353A_0r0[31:0], L353A_0r1[31:0], L353A_0a, L199_0r0[31:0], L199_0r1[31:0], L199_0a, L345A_0r0, L345A_0r1, L345A_0a, reset);
  tkf32mo0w0_o0w32 I84 (L264P_0r0[31:0], L264P_0r1[31:0], L264P_0a, L320A_0r, L320A_0a, L321_0r0[31:0], L321_0r1[31:0], L321_0a, reset);
  tkf32mo0w0_o0w32 I85 (L8_0r0[31:0], L8_0r1[31:0], L8_0a, L322_0r, L322_0a, L323_0r0[31:0], L323_0r1[31:0], L323_0a, reset);
  tkm2x32b I86 (L321_0r0[31:0], L321_0r1[31:0], L321_0a, L323_0r0[31:0], L323_0r1[31:0], L323_0a, L318A_0r0[31:0], L318A_0r1[31:0], L318A_0a, reset);
  tko0m2_1nm2b1 I87 (L320P_0r, L320P_0a, L324A_0r0[1:0], L324A_0r1[1:0], L324A_0a, reset);
  tko0m2_1nm2b2 I88 (L322_0r, L322_0a, L325_0r0[1:0], L325_0r1[1:0], L325_0a, reset);
  tkm2x2b I89 (L324P_0r0[1:0], L324P_0r1[1:0], L324P_0a, L325_0r0[1:0], L325_0r1[1:0], L325_0a, L326A_0r0[1:0], L326A_0r1[1:0], L326A_0a, reset);
  tkj2m0_2 I90 (L319P_0r, L319P_0a, L326P_0r0[1:0], L326P_0r1[1:0], L326P_0a, L327A_0r0[1:0], L327A_0r1[1:0], L327A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I91 (L327P_0r0[1:0], L327P_0r1[1:0], L327P_0a, L267_0r, L267_0a, L9_0r, L9_0a, reset);
  tkvaV32_wo0w32_ro0w32o0w32 I92 (L318P_0r0[31:0], L318P_0r1[31:0], L318P_0a, L319A_0r, L319A_0a, L367P_0r, L367P_0a, L385P_0r, L385P_0a, a_0r0[31:0], a_0r1[31:0], a_0a, L169_0r0[31:0], L169_0r1[31:0], L169_0a, reset);
  tkj32m32_0 I93 (x_0r0[31:0], x_0r1[31:0], x_0a, L284P_0r, L284P_0a, L4A_0r0[31:0], L4A_0r1[31:0], L4A_0a, reset);
  tko0m2_1nm2b1 I94 (L7_0r, L7_0a, L332_0r0[1:0], L332_0r1[1:0], L332_0a, reset);
  tko0m2_1nm2b2 I95 (L253P_0r, L253P_0a, L333A_0r0[1:0], L333A_0r1[1:0], L333A_0a, reset);
  tkm2x2b I96 (L332_0r0[1:0], L332_0r1[1:0], L332_0a, L333P_0r0[1:0], L333P_0r1[1:0], L333P_0a, L334A_0r0[1:0], L334A_0r1[1:0], L334A_0a, reset);
  tkj34m32_2 I97 (coefs_2_0r0[31:0], coefs_2_0r1[31:0], coefs_2_0a, L334P_0r0[1:0], L334P_0r1[1:0], L334P_0a, L335_0r0[33:0], L335_0r1[33:0], L335_0a, reset);
  tks34_o32w2_1o0w32_2o0w32 I98 (L335_0r0[33:0], L335_0r1[33:0], L335_0a, L8_0r0[31:0], L8_0r1[31:0], L8_0a, L249_0r0[31:0], L249_0r1[31:0], L249_0a, reset);
  tki I99 (L281P_0r, L281P_0a, L284A_0r, L284A_0a, reset);
  tkj64m32_32_0 I100 (L211_0r0[31:0], L211_0r1[31:0], L211_0a, coefs_0_0r0[31:0], coefs_0_0r1[31:0], coefs_0_0a, L217_0r, L217_0a, L206_0r0[63:0], L206_0r1[63:0], L206_0a, reset);
  tkj64m32_32_0 I101 (L229_0r0[31:0], L229_0r1[31:0], L229_0a, coefs_1_0r0[31:0], coefs_1_0r1[31:0], coefs_1_0a, L235_0r, L235_0a, L224_0r0[63:0], L224_0r1[63:0], L224_0a, reset);
  tkj64m32_32 I102 (L247_0r0[31:0], L247_0r1[31:0], L247_0a, L249_0r0[31:0], L249_0r1[31:0], L249_0a, L242_0r0[63:0], L242_0r1[63:0], L242_0a, reset);
  tko1m1_1nm1b1_2nei0w1bt1o0w1b I103 (L345P_0r0, L345P_0r1, L345P_0a, L21_0r0, L21_0r1, L21_0a, reset);
  tko1m1_1nm1b1_2eqi0w1bt1o0w1b I104 (L346P_0r0, L346P_0r1, L346P_0a, L54_0r0, L54_0r1, L54_0a, reset);
  tko3m4_1nm1b0_2api0w3bt1o0w1b_3nm4b1_4addt2o0w4bt3o0w4b I105 (L347P_0r0[2:0], L347P_0r1[2:0], L347P_0a, L68_0r0[3:0], L68_0r1[3:0], L68_0a, reset);
  tko1m1_1nm1b1_2eqi0w1bt1o0w1b I106 (L348P_0r0, L348P_0r1, L348P_0a, L80_0r0, L80_0r1, L80_0a, reset);
  tko3m4_1nm1b0_2api0w3bt1o0w1b_3nm4b1_4addt2o0w4bt3o0w4b I107 (L349_0r0[2:0], L349_0r1[2:0], L349_0a, L94A_0r0[3:0], L94A_0r1[3:0], L94A_0a, reset);
  tko32m1_1nm32b0_2sgti0w32bt1o0w32b I108 (L350_0r0[31:0], L350_0r1[31:0], L350_0a, L106_0r0, L106_0r1, L106_0a, reset);
  tko32m33_1api0w32bi31w1b_2nm33b1_3subt1o0w33bt2o0w33b I109 (L351_0r0[31:0], L351_0r1[31:0], L351_0a, L125A_0r0[32:0], L125A_0r1[32:0], L125A_0a, reset);
  tko3m1_1nm3b1_2eqi0w3bt1o0w3b I110 (L352_0r0[2:0], L352_0r1[2:0], L352_0a, L136_0r0, L136_0r1, L136_0a, reset);
  tko32m33_1api0w32bi31w1b_2nm33b1_3subt1o0w33bt2o0w33b I111 (L353P_0r0[31:0], L353P_0r1[31:0], L353P_0a, L272A_0r0[32:0], L272A_0r1[32:0], L272A_0a, reset);
  tkj32m32_0_0_0 I112 (L302P_0r0[31:0], L302P_0r1[31:0], L302P_0a, L257P_0r, L257P_0a, L148P_0r, L148P_0a, L255P_0r, L255P_0a, L264A_0r0[31:0], L264A_0r1[31:0], L264A_0a, reset);
  tkf0mo0w0_o0w0 I113 (L140_0r, L140_0a, L363A_0r, L363A_0a, L187A_0r, L187A_0a, reset);
  tkf0mo0w0_o0w0 I114 (L145P_0r, L145P_0a, L366A_0r, L366A_0a, L148A_0r, L148A_0a, reset);
  tkf0mo0w0_o0w0 I115 (L278_0r, L278_0a, L367A_0r, L367A_0a, L281A_0r, L281A_0a, reset);
  tkm3x32b I116 (L299_0r0[31:0], L299_0r1[31:0], L299_0a, L295_0r0[31:0], L295_0r1[31:0], L295_0a, L297_0r0[31:0], L297_0r1[31:0], L297_0a, L395A_0r0[31:0], L395A_0r1[31:0], L395A_0a, reset);
  tkf32mo0w0_o0w32 I117 (L395P_0r0[31:0], L395P_0r1[31:0], L395P_0a, L338A_0r, L338A_0a, L302A_0r0[31:0], L302A_0r1[31:0], L302A_0a, reset);
  tko64m32_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b_4apt3o0w32b I118 (L206_0r0[63:0], L206_0r1[63:0], L206_0a, L295_0r0[31:0], L295_0r1[31:0], L295_0a, reset);
  tko64m32_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b_4apt3o0w32b I119 (L224_0r0[63:0], L224_0r1[63:0], L224_0a, L297_0r0[31:0], L297_0r1[31:0], L297_0a, reset);
  tko64m32_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b_4apt3o0w32b I120 (L242_0r0[63:0], L242_0r1[63:0], L242_0a, L299_0r0[31:0], L299_0r1[31:0], L299_0a, reset);
  tkl32x1 I121 (L4A_0r0[31:0], L4A_0r1[31:0], L4A_0a, L4P_0r0[31:0], L4P_0r1[31:0], L4P_0a, reset);
  tkl0x1 I122 (L13A_0r, L13A_0a, L13P_0r, L13P_0a, reset);
  tkl0x1 I123 (L14A_0r, L14A_0a, L14P_0r, L14P_0a, reset);
  tkl0x1 I124 (L16A_0r, L16A_0a, L16P_0r, L16P_0a, reset);
  tkl0x1 I125 (L49A_0r, L49A_0a, L49P_0r, L49P_0a, reset);
  tkl0x1 I126 (L56A_0r, L56A_0a, L56P_0r, L56P_0a, reset);
  tkl0x1 I127 (L63A_0r, L63A_0a, L63P_0r, L63P_0a, reset);
  tkl0x1 I128 (L72A_0r, L72A_0a, L72P_0r, L72P_0a, reset);
  tkl0x1 I129 (L73A_0r, L73A_0a, L73P_0r, L73P_0a, reset);
  tkl0x1 I130 (L75A_0r, L75A_0a, L75P_0r, L75P_0a, reset);
  tkl0x1 I131 (L82A_0r, L82A_0a, L82P_0r, L82P_0a, reset);
  tkl0x1 I132 (L89A_0r, L89A_0a, L89P_0r, L89P_0a, reset);
  tkl4x1 I133 (L94A_0r0[3:0], L94A_0r1[3:0], L94A_0a, L94P_0r0[3:0], L94P_0r1[3:0], L94P_0a, reset);
  tkl0x1 I134 (L98A_0r, L98A_0a, L98P_0r, L98P_0a, reset);
  tkl0x1 I135 (L99A_0r, L99A_0a, L99P_0r, L99P_0a, reset);
  tkl0x1 I136 (L101A_0r, L101A_0a, L101P_0r, L101P_0a, reset);
  tkl0x1 I137 (L110A_0r, L110A_0a, L110P_0r, L110P_0a, reset);
  tkl32x1 I138 (L111A_0r0[31:0], L111A_0r1[31:0], L111A_0a, L111P_0r0[31:0], L111P_0r1[31:0], L111P_0a, reset);
  tkl0x1 I139 (L112A_0r, L112A_0a, L112P_0r, L112P_0a, reset);
  tkl64x1 I140 (L114A_0r0[63:0], L114A_0r1[63:0], L114A_0a, L114P_0r0[63:0], L114P_0r1[63:0], L114P_0a, reset);
  tkl0x1 I141 (L116A_0r, L116A_0a, L116P_0r, L116P_0a, reset);
  tkl0x1 I142 (L120A_0r, L120A_0a, L120P_0r, L120P_0a, reset);
  tkl33x1 I143 (L125A_0r0[32:0], L125A_0r1[32:0], L125A_0a, L125P_0r0[32:0], L125P_0r1[32:0], L125P_0a, reset);
  tkl0x1 I144 (L128A_0r, L128A_0a, L128P_0r, L128P_0a, reset);
  tkl0x1 I145 (L131A_0r, L131A_0a, L131P_0r, L131P_0a, reset);
  tkl0x1 I146 (L145A_0r, L145A_0a, L145P_0r, L145P_0a, reset);
  tkl0x1 I147 (L148A_0r, L148A_0a, L148P_0r, L148P_0a, reset);
  tkl3x1 I148 (L149A_0r0[2:0], L149A_0r1[2:0], L149A_0a, L149P_0r0[2:0], L149P_0r1[2:0], L149P_0a, reset);
  tkl0x1 I149 (L150A_0r, L150A_0a, L150P_0r, L150P_0a, reset);
  tkl0x1 I150 (L151A_0r, L151A_0a, L151P_0r, L151P_0a, reset);
  tkl3x1 I151 (L152A_0r0[2:0], L152A_0r1[2:0], L152A_0a, L152P_0r0[2:0], L152P_0r1[2:0], L152P_0a, reset);
  tkl0x1 I152 (L153A_0r, L153A_0a, L153P_0r, L153P_0a, reset);
  tkl3x1 I153 (L154A_0r0[2:0], L154A_0r1[2:0], L154A_0a, L154P_0r0[2:0], L154P_0r1[2:0], L154P_0a, reset);
  tkl3x1 I154 (L156A_0r0[2:0], L156A_0r1[2:0], L156A_0a, L156P_0r0[2:0], L156P_0r1[2:0], L156P_0a, reset);
  tkl3x1 I155 (L157A_0r0[2:0], L157A_0r1[2:0], L157A_0a, L157P_0r0[2:0], L157P_0r1[2:0], L157P_0a, reset);
  tkl3x1 I156 (L158A_0r0[2:0], L158A_0r1[2:0], L158A_0a, L158P_0r0[2:0], L158P_0r1[2:0], L158P_0a, reset);
  tkl3x1 I157 (L160A_0r0[2:0], L160A_0r1[2:0], L160A_0a, L160P_0r0[2:0], L160P_0r1[2:0], L160P_0a, reset);
  tkl3x1 I158 (L161A_0r0[2:0], L161A_0r1[2:0], L161A_0a, L161P_0r0[2:0], L161P_0r1[2:0], L161P_0a, reset);
  tkl32x1 I159 (L162A_0r0[31:0], L162A_0r1[31:0], L162A_0a, L162P_0r0[31:0], L162P_0r1[31:0], L162P_0a, reset);
  tkl0x1 I160 (L163A_0r, L163A_0a, L163P_0r, L163P_0a, reset);
  tkl32x1 I161 (L165A_0r0[31:0], L165A_0r1[31:0], L165A_0a, L165P_0r0[31:0], L165P_0r1[31:0], L165P_0a, reset);
  tkl32x1 I162 (L167A_0r0[31:0], L167A_0r1[31:0], L167A_0a, L167P_0r0[31:0], L167P_0r1[31:0], L167P_0a, reset);
  tkl3x1 I163 (L170A_0r0[2:0], L170A_0r1[2:0], L170A_0a, L170P_0r0[2:0], L170P_0r1[2:0], L170P_0a, reset);
  tkl3x1 I164 (L171A_0r0[2:0], L171A_0r1[2:0], L171A_0a, L171P_0r0[2:0], L171P_0r1[2:0], L171P_0a, reset);
  tkl3x1 I165 (L172A_0r0[2:0], L172A_0r1[2:0], L172A_0a, L172P_0r0[2:0], L172P_0r1[2:0], L172P_0a, reset);
  tkl3x1 I166 (L173A_0r0[2:0], L173A_0r1[2:0], L173A_0a, L173P_0r0[2:0], L173P_0r1[2:0], L173P_0a, reset);
  tkl3x1 I167 (L174A_0r0[2:0], L174A_0r1[2:0], L174A_0a, L174P_0r0[2:0], L174P_0r1[2:0], L174P_0a, reset);
  tkl32x1 I168 (L175A_0r0[31:0], L175A_0r1[31:0], L175A_0a, L175P_0r0[31:0], L175P_0r1[31:0], L175P_0a, reset);
  tkl0x1 I169 (L176A_0r, L176A_0a, L176P_0r, L176P_0a, reset);
  tkl0x1 I170 (L177A_0r, L177A_0a, L177P_0r, L177P_0a, reset);
  tkl32x1 I171 (L178A_0r0[31:0], L178A_0r1[31:0], L178A_0a, L178P_0r0[31:0], L178P_0r1[31:0], L178P_0a, reset);
  tkl32x1 I172 (L180A_0r0[31:0], L180A_0r1[31:0], L180A_0a, L180P_0r0[31:0], L180P_0r1[31:0], L180P_0a, reset);
  tkl2x1 I173 (L181A_0r0[1:0], L181A_0r1[1:0], L181A_0a, L181P_0r0[1:0], L181P_0r1[1:0], L181P_0a, reset);
  tkl2x1 I174 (L183A_0r0[1:0], L183A_0r1[1:0], L183A_0a, L183P_0r0[1:0], L183P_0r1[1:0], L183P_0a, reset);
  tkl2x1 I175 (L184A_0r0[1:0], L184A_0r1[1:0], L184A_0a, L184P_0r0[1:0], L184P_0r1[1:0], L184P_0a, reset);
  tkl32x1 I176 (L185A_0r0[31:0], L185A_0r1[31:0], L185A_0a, L185P_0r0[31:0], L185P_0r1[31:0], L185P_0a, reset);
  tkl0x1 I177 (L186A_0r, L186A_0a, L186P_0r, L186P_0a, reset);
  tkl0x1 I178 (L187A_0r, L187A_0a, L187P_0r, L187P_0a, reset);
  tkl32x1 I179 (L188A_0r0[31:0], L188A_0r1[31:0], L188A_0a, L188P_0r0[31:0], L188P_0r1[31:0], L188P_0a, reset);
  tkl0x1 I180 (L189A_0r, L189A_0a, L189P_0r, L189P_0a, reset);
  tkl3x1 I181 (L193A_0r0[2:0], L193A_0r1[2:0], L193A_0a, L193P_0r0[2:0], L193P_0r1[2:0], L193P_0a, reset);
  tkl3x1 I182 (L194A_0r0[2:0], L194A_0r1[2:0], L194A_0a, L194P_0r0[2:0], L194P_0r1[2:0], L194P_0a, reset);
  tkl3x1 I183 (L196A_0r0[2:0], L196A_0r1[2:0], L196A_0a, L196P_0r0[2:0], L196P_0r1[2:0], L196P_0a, reset);
  tkl3x1 I184 (L197A_0r0[2:0], L197A_0r1[2:0], L197A_0a, L197P_0r0[2:0], L197P_0r1[2:0], L197P_0a, reset);
  tkl0x1 I185 (L198A_0r, L198A_0a, L198P_0r, L198P_0a, reset);
  tkl0x1 I186 (L253A_0r, L253A_0a, L253P_0r, L253P_0a, reset);
  tkl0x1 I187 (L255A_0r, L255A_0a, L255P_0r, L255P_0a, reset);
  tkl0x1 I188 (L257A_0r, L257A_0a, L257P_0r, L257P_0a, reset);
  tkl0x1 I189 (L260A_0r, L260A_0a, L260P_0r, L260P_0a, reset);
  tkl32x1 I190 (L264A_0r0[31:0], L264A_0r1[31:0], L264A_0a, L264P_0r0[31:0], L264P_0r1[31:0], L264P_0a, reset);
  tkl33x1 I191 (L272A_0r0[32:0], L272A_0r1[32:0], L272A_0a, L272P_0r0[32:0], L272P_0r1[32:0], L272P_0a, reset);
  tkl0x1 I192 (L275A_0r, L275A_0a, L275P_0r, L275P_0a, reset);
  tkl0x1 I193 (L277A_0r, L277A_0a, L277P_0r, L277P_0a, reset);
  tkl0x1 I194 (L281A_0r, L281A_0a, L281P_0r, L281P_0a, reset);
  tkl0x1 I195 (L284A_0r, L284A_0a, L284P_0r, L284P_0a, reset);
  tkl32x1 I196 (L302A_0r0[31:0], L302A_0r1[31:0], L302A_0a, L302P_0r0[31:0], L302P_0r1[31:0], L302P_0a, reset);
  tkl32x1 I197 (L308A_0r0[31:0], L308A_0r1[31:0], L308A_0a, L308P_0r0[31:0], L308P_0r1[31:0], L308P_0a, reset);
  tkl32x1 I198 (L313A_0r0[31:0], L313A_0r1[31:0], L313A_0a, L313P_0r0[31:0], L313P_0r1[31:0], L313P_0a, reset);
  tkl2x1 I199 (L317A_0r0[1:0], L317A_0r1[1:0], L317A_0a, L317P_0r0[1:0], L317P_0r1[1:0], L317P_0a, reset);
  tkl32x1 I200 (L318A_0r0[31:0], L318A_0r1[31:0], L318A_0a, L318P_0r0[31:0], L318P_0r1[31:0], L318P_0a, reset);
  tkl0x1 I201 (L319A_0r, L319A_0a, L319P_0r, L319P_0a, reset);
  tkl0x1 I202 (L320A_0r, L320A_0a, L320P_0r, L320P_0a, reset);
  tkl2x1 I203 (L324A_0r0[1:0], L324A_0r1[1:0], L324A_0a, L324P_0r0[1:0], L324P_0r1[1:0], L324P_0a, reset);
  tkl2x1 I204 (L326A_0r0[1:0], L326A_0r1[1:0], L326A_0a, L326P_0r0[1:0], L326P_0r1[1:0], L326P_0a, reset);
  tkl2x1 I205 (L327A_0r0[1:0], L327A_0r1[1:0], L327A_0a, L327P_0r0[1:0], L327P_0r1[1:0], L327P_0a, reset);
  tkl2x1 I206 (L333A_0r0[1:0], L333A_0r1[1:0], L333A_0a, L333P_0r0[1:0], L333P_0r1[1:0], L333P_0a, reset);
  tkl2x1 I207 (L334A_0r0[1:0], L334A_0r1[1:0], L334A_0a, L334P_0r0[1:0], L334P_0r1[1:0], L334P_0a, reset);
  tkl0x1 I208 (L338A_0r, L338A_0a, L338P_0r, L338P_0a, reset);
  tkl1x1 I209 (L345A_0r0, L345A_0r1, L345A_0a, L345P_0r0, L345P_0r1, L345P_0a, reset);
  tkl1x1 I210 (L346A_0r0, L346A_0r1, L346A_0a, L346P_0r0, L346P_0r1, L346P_0a, reset);
  tkl3x1 I211 (L347A_0r0[2:0], L347A_0r1[2:0], L347A_0a, L347P_0r0[2:0], L347P_0r1[2:0], L347P_0a, reset);
  tkl1x1 I212 (L348A_0r0, L348A_0r1, L348A_0a, L348P_0r0, L348P_0r1, L348P_0a, reset);
  tkl32x1 I213 (L353A_0r0[31:0], L353A_0r1[31:0], L353A_0a, L353P_0r0[31:0], L353P_0r1[31:0], L353P_0a, reset);
  tkl32x1 I214 (L358A_0r0[31:0], L358A_0r1[31:0], L358A_0a, L358P_0r0[31:0], L358P_0r1[31:0], L358P_0a, reset);
  tkl32x1 I215 (L359A_0r0[31:0], L359A_0r1[31:0], L359A_0a, L359P_0r0[31:0], L359P_0r1[31:0], L359P_0a, reset);
  tkl32x1 I216 (L360A_0r0[31:0], L360A_0r1[31:0], L360A_0a, L360P_0r0[31:0], L360P_0r1[31:0], L360P_0a, reset);
  tkl0x1 I217 (L361A_0r, L361A_0a, L361P_0r, L361P_0a, reset);
  tkl0x1 I218 (L362A_0r, L362A_0a, L362P_0r, L362P_0a, reset);
  tkl0x1 I219 (L363A_0r, L363A_0a, L363P_0r, L363P_0a, reset);
  tkl0x1 I220 (L364A_0r, L364A_0a, L364P_0r, L364P_0a, reset);
  tkl0x1 I221 (L366A_0r, L366A_0a, L366P_0r, L366P_0a, reset);
  tkl0x1 I222 (L367A_0r, L367A_0a, L367P_0r, L367P_0a, reset);
  tkl0x1 I223 (L385A_0r, L385A_0a, L385P_0r, L385P_0a, reset);
  tkl32x1 I224 (L395A_0r0[31:0], L395A_0r1[31:0], L395A_0a, L395P_0r0[31:0], L395P_0r1[31:0], L395P_0a, reset);
  tkr_dr_monitor #("Poly_eval.L4.P", 32) I225 (L4P_0r0[31:0], L4P_0r1[31:0], L4P_0a);
  tkr_dr_monitor #("Poly_eval.L4.A", 32) I226 (L4A_0r0[31:0], L4A_0r1[31:0], L4A_0a);
  tkr_ra_monitor #("Poly_eval.L7.L") I227 (L7_0r, L7_0a);
  tkr_dr_monitor #("Poly_eval.L8.L", 32) I228 (L8_0r0[31:0], L8_0r1[31:0], L8_0a);
  tkr_ra_monitor #("Poly_eval.L9.L") I229 (L9_0r, L9_0a);
  tkr_ra_monitor #("Poly_eval.L13.P") I230 (L13P_0r, L13P_0a);
  tkr_ra_monitor #("Poly_eval.L13.A") I231 (L13A_0r, L13A_0a);
  tkr_ra_monitor #("Poly_eval.L14.P") I232 (L14P_0r, L14P_0a);
  tkr_ra_monitor #("Poly_eval.L14.A") I233 (L14A_0r, L14A_0a);
  tkr_ra_monitor #("Poly_eval.L16.P") I234 (L16P_0r, L16P_0a);
  tkr_ra_monitor #("Poly_eval.L16.A") I235 (L16A_0r, L16A_0a);
  tkr_dr_monitor #("Poly_eval.L21.L", 1) I236 (L21_0r0, L21_0r1, L21_0a);
  tkr_ra_monitor #("Poly_eval.L38.L") I237 (L38_0r, L38_0a);
  tkr_dr_monitor #("Poly_eval.L39.L", 32) I238 (L39_0r0[31:0], L39_0r1[31:0], L39_0a);
  tkr_ra_monitor #("Poly_eval.L41.L") I239 (L41_0r, L41_0a);
  tkr_ra_monitor #("Poly_eval.L45.L") I240 (L45_0r, L45_0a);
  tkr_ra_monitor #("Poly_eval.L49.P") I241 (L49P_0r, L49P_0a);
  tkr_ra_monitor #("Poly_eval.L49.A") I242 (L49A_0r, L49A_0a);
  tkr_dr_monitor #("Poly_eval.L54.L", 1) I243 (L54_0r0, L54_0r1, L54_0a);
  tkr_ra_monitor #("Poly_eval.L56.P") I244 (L56P_0r, L56P_0a);
  tkr_ra_monitor #("Poly_eval.L56.A") I245 (L56A_0r, L56A_0a);
  tkr_ra_monitor #("Poly_eval.L61.L") I246 (L61_0r, L61_0a);
  tkr_ra_monitor #("Poly_eval.L63.P") I247 (L63P_0r, L63P_0a);
  tkr_ra_monitor #("Poly_eval.L63.A") I248 (L63A_0r, L63A_0a);
  tkr_dr_monitor #("Poly_eval.L68.L", 4) I249 (L68_0r0[3:0], L68_0r1[3:0], L68_0a);
  tkr_ra_monitor #("Poly_eval.L71.L") I250 (L71_0r, L71_0a);
  tkr_ra_monitor #("Poly_eval.L72.P") I251 (L72P_0r, L72P_0a);
  tkr_ra_monitor #("Poly_eval.L72.A") I252 (L72A_0r, L72A_0a);
  tkr_ra_monitor #("Poly_eval.L73.P") I253 (L73P_0r, L73P_0a);
  tkr_ra_monitor #("Poly_eval.L73.A") I254 (L73A_0r, L73A_0a);
  tkr_ra_monitor #("Poly_eval.L75.P") I255 (L75P_0r, L75P_0a);
  tkr_ra_monitor #("Poly_eval.L75.A") I256 (L75A_0r, L75A_0a);
  tkr_dr_monitor #("Poly_eval.L80.L", 1) I257 (L80_0r0, L80_0r1, L80_0a);
  tkr_ra_monitor #("Poly_eval.L82.P") I258 (L82P_0r, L82P_0a);
  tkr_ra_monitor #("Poly_eval.L82.A") I259 (L82A_0r, L82A_0a);
  tkr_ra_monitor #("Poly_eval.L87.L") I260 (L87_0r, L87_0a);
  tkr_ra_monitor #("Poly_eval.L89.P") I261 (L89P_0r, L89P_0a);
  tkr_ra_monitor #("Poly_eval.L89.A") I262 (L89A_0r, L89A_0a);
  tkr_dr_monitor #("Poly_eval.L94.P", 4) I263 (L94P_0r0[3:0], L94P_0r1[3:0], L94P_0a);
  tkr_dr_monitor #("Poly_eval.L94.A", 4) I264 (L94A_0r0[3:0], L94A_0r1[3:0], L94A_0a);
  tkr_ra_monitor #("Poly_eval.L97.L") I265 (L97_0r, L97_0a);
  tkr_ra_monitor #("Poly_eval.L98.P") I266 (L98P_0r, L98P_0a);
  tkr_ra_monitor #("Poly_eval.L98.A") I267 (L98A_0r, L98A_0a);
  tkr_ra_monitor #("Poly_eval.L99.P") I268 (L99P_0r, L99P_0a);
  tkr_ra_monitor #("Poly_eval.L99.A") I269 (L99A_0r, L99A_0a);
  tkr_ra_monitor #("Poly_eval.L101.P") I270 (L101P_0r, L101P_0a);
  tkr_ra_monitor #("Poly_eval.L101.A") I271 (L101A_0r, L101A_0a);
  tkr_dr_monitor #("Poly_eval.L106.L", 1) I272 (L106_0r0, L106_0r1, L106_0a);
  tkr_ra_monitor #("Poly_eval.L110.P") I273 (L110P_0r, L110P_0a);
  tkr_ra_monitor #("Poly_eval.L110.A") I274 (L110A_0r, L110A_0a);
  tkr_dr_monitor #("Poly_eval.L111.P", 32) I275 (L111P_0r0[31:0], L111P_0r1[31:0], L111P_0a);
  tkr_dr_monitor #("Poly_eval.L111.A", 32) I276 (L111A_0r0[31:0], L111A_0r1[31:0], L111A_0a);
  tkr_ra_monitor #("Poly_eval.L112.P") I277 (L112P_0r, L112P_0a);
  tkr_ra_monitor #("Poly_eval.L112.A") I278 (L112A_0r, L112A_0a);
  tkr_dr_monitor #("Poly_eval.L113.L", 32) I279 (L113_0r0[31:0], L113_0r1[31:0], L113_0a);
  tkr_dr_monitor #("Poly_eval.L114.P", 64) I280 (L114P_0r0[63:0], L114P_0r1[63:0], L114P_0a);
  tkr_dr_monitor #("Poly_eval.L114.A", 64) I281 (L114A_0r0[63:0], L114A_0r1[63:0], L114A_0a);
  tkr_dr_monitor #("Poly_eval.L115.L", 33) I282 (L115_0r0[32:0], L115_0r1[32:0], L115_0a);
  tkr_ra_monitor #("Poly_eval.L116.P") I283 (L116P_0r, L116P_0a);
  tkr_ra_monitor #("Poly_eval.L116.A") I284 (L116A_0r, L116A_0a);
  tkr_ra_monitor #("Poly_eval.L120.P") I285 (L120P_0r, L120P_0a);
  tkr_ra_monitor #("Poly_eval.L120.A") I286 (L120A_0r, L120A_0a);
  tkr_dr_monitor #("Poly_eval.L125.P", 33) I287 (L125P_0r0[32:0], L125P_0r1[32:0], L125P_0a);
  tkr_dr_monitor #("Poly_eval.L125.A", 33) I288 (L125A_0r0[32:0], L125A_0r1[32:0], L125A_0a);
  tkr_ra_monitor #("Poly_eval.L128.P") I289 (L128P_0r, L128P_0a);
  tkr_ra_monitor #("Poly_eval.L128.A") I290 (L128A_0r, L128A_0a);
  tkr_ra_monitor #("Poly_eval.L131.P") I291 (L131P_0r, L131P_0a);
  tkr_ra_monitor #("Poly_eval.L131.A") I292 (L131A_0r, L131A_0a);
  tkr_dr_monitor #("Poly_eval.L136.L", 1) I293 (L136_0r0, L136_0r1, L136_0a);
  tkr_ra_monitor #("Poly_eval.L138.L") I294 (L138_0r, L138_0a);
  tkr_ra_monitor #("Poly_eval.L140.L") I295 (L140_0r, L140_0a);
  tkr_ra_monitor #("Poly_eval.L143.L") I296 (L143_0r, L143_0a);
  tkr_ra_monitor #("Poly_eval.L145.P") I297 (L145P_0r, L145P_0a);
  tkr_ra_monitor #("Poly_eval.L145.A") I298 (L145A_0r, L145A_0a);
  tkr_ra_monitor #("Poly_eval.L148.P") I299 (L148P_0r, L148P_0a);
  tkr_ra_monitor #("Poly_eval.L148.A") I300 (L148A_0r, L148A_0a);
  tkr_dr_monitor #("Poly_eval.L149.P", 3) I301 (L149P_0r0[2:0], L149P_0r1[2:0], L149P_0a);
  tkr_dr_monitor #("Poly_eval.L149.A", 3) I302 (L149A_0r0[2:0], L149A_0r1[2:0], L149A_0a);
  tkr_ra_monitor #("Poly_eval.L150.P") I303 (L150P_0r, L150P_0a);
  tkr_ra_monitor #("Poly_eval.L150.A") I304 (L150A_0r, L150A_0a);
  tkr_ra_monitor #("Poly_eval.L151.P") I305 (L151P_0r, L151P_0a);
  tkr_ra_monitor #("Poly_eval.L151.A") I306 (L151A_0r, L151A_0a);
  tkr_dr_monitor #("Poly_eval.L152.P", 3) I307 (L152P_0r0[2:0], L152P_0r1[2:0], L152P_0a);
  tkr_dr_monitor #("Poly_eval.L152.A", 3) I308 (L152A_0r0[2:0], L152A_0r1[2:0], L152A_0a);
  tkr_ra_monitor #("Poly_eval.L153.P") I309 (L153P_0r, L153P_0a);
  tkr_ra_monitor #("Poly_eval.L153.A") I310 (L153A_0r, L153A_0a);
  tkr_dr_monitor #("Poly_eval.L154.P", 3) I311 (L154P_0r0[2:0], L154P_0r1[2:0], L154P_0a);
  tkr_dr_monitor #("Poly_eval.L154.A", 3) I312 (L154A_0r0[2:0], L154A_0r1[2:0], L154A_0a);
  tkr_ra_monitor #("Poly_eval.L155.L") I313 (L155_0r, L155_0a);
  tkr_dr_monitor #("Poly_eval.L156.P", 3) I314 (L156P_0r0[2:0], L156P_0r1[2:0], L156P_0a);
  tkr_dr_monitor #("Poly_eval.L156.A", 3) I315 (L156A_0r0[2:0], L156A_0r1[2:0], L156A_0a);
  tkr_dr_monitor #("Poly_eval.L157.P", 3) I316 (L157P_0r0[2:0], L157P_0r1[2:0], L157P_0a);
  tkr_dr_monitor #("Poly_eval.L157.A", 3) I317 (L157A_0r0[2:0], L157A_0r1[2:0], L157A_0a);
  tkr_dr_monitor #("Poly_eval.L158.P", 3) I318 (L158P_0r0[2:0], L158P_0r1[2:0], L158P_0a);
  tkr_dr_monitor #("Poly_eval.L158.A", 3) I319 (L158A_0r0[2:0], L158A_0r1[2:0], L158A_0a);
  tkr_dr_monitor #("Poly_eval.L159.L", 3) I320 (L159_0r0[2:0], L159_0r1[2:0], L159_0a);
  tkr_dr_monitor #("Poly_eval.L160.P", 3) I321 (L160P_0r0[2:0], L160P_0r1[2:0], L160P_0a);
  tkr_dr_monitor #("Poly_eval.L160.A", 3) I322 (L160A_0r0[2:0], L160A_0r1[2:0], L160A_0a);
  tkr_dr_monitor #("Poly_eval.L161.P", 3) I323 (L161P_0r0[2:0], L161P_0r1[2:0], L161P_0a);
  tkr_dr_monitor #("Poly_eval.L161.A", 3) I324 (L161A_0r0[2:0], L161A_0r1[2:0], L161A_0a);
  tkr_dr_monitor #("Poly_eval.L162.P", 32) I325 (L162P_0r0[31:0], L162P_0r1[31:0], L162P_0a);
  tkr_dr_monitor #("Poly_eval.L162.A", 32) I326 (L162A_0r0[31:0], L162A_0r1[31:0], L162A_0a);
  tkr_ra_monitor #("Poly_eval.L163.P") I327 (L163P_0r, L163P_0a);
  tkr_ra_monitor #("Poly_eval.L163.A") I328 (L163A_0r, L163A_0a);
  tkr_ra_monitor #("Poly_eval.L164.L") I329 (L164_0r, L164_0a);
  tkr_dr_monitor #("Poly_eval.L165.P", 32) I330 (L165P_0r0[31:0], L165P_0r1[31:0], L165P_0a);
  tkr_dr_monitor #("Poly_eval.L165.A", 32) I331 (L165A_0r0[31:0], L165A_0r1[31:0], L165A_0a);
  tkr_ra_monitor #("Poly_eval.L166.L") I332 (L166_0r, L166_0a);
  tkr_dr_monitor #("Poly_eval.L167.P", 32) I333 (L167P_0r0[31:0], L167P_0r1[31:0], L167P_0a);
  tkr_dr_monitor #("Poly_eval.L167.A", 32) I334 (L167A_0r0[31:0], L167A_0r1[31:0], L167A_0a);
  tkr_ra_monitor #("Poly_eval.L168.L") I335 (L168_0r, L168_0a);
  tkr_dr_monitor #("Poly_eval.L169.L", 32) I336 (L169_0r0[31:0], L169_0r1[31:0], L169_0a);
  tkr_dr_monitor #("Poly_eval.L170.P", 3) I337 (L170P_0r0[2:0], L170P_0r1[2:0], L170P_0a);
  tkr_dr_monitor #("Poly_eval.L170.A", 3) I338 (L170A_0r0[2:0], L170A_0r1[2:0], L170A_0a);
  tkr_dr_monitor #("Poly_eval.L171.P", 3) I339 (L171P_0r0[2:0], L171P_0r1[2:0], L171P_0a);
  tkr_dr_monitor #("Poly_eval.L171.A", 3) I340 (L171A_0r0[2:0], L171A_0r1[2:0], L171A_0a);
  tkr_dr_monitor #("Poly_eval.L172.P", 3) I341 (L172P_0r0[2:0], L172P_0r1[2:0], L172P_0a);
  tkr_dr_monitor #("Poly_eval.L172.A", 3) I342 (L172A_0r0[2:0], L172A_0r1[2:0], L172A_0a);
  tkr_dr_monitor #("Poly_eval.L173.P", 3) I343 (L173P_0r0[2:0], L173P_0r1[2:0], L173P_0a);
  tkr_dr_monitor #("Poly_eval.L173.A", 3) I344 (L173A_0r0[2:0], L173A_0r1[2:0], L173A_0a);
  tkr_dr_monitor #("Poly_eval.L174.P", 3) I345 (L174P_0r0[2:0], L174P_0r1[2:0], L174P_0a);
  tkr_dr_monitor #("Poly_eval.L174.A", 3) I346 (L174A_0r0[2:0], L174A_0r1[2:0], L174A_0a);
  tkr_dr_monitor #("Poly_eval.L175.P", 32) I347 (L175P_0r0[31:0], L175P_0r1[31:0], L175P_0a);
  tkr_dr_monitor #("Poly_eval.L175.A", 32) I348 (L175A_0r0[31:0], L175A_0r1[31:0], L175A_0a);
  tkr_ra_monitor #("Poly_eval.L176.P") I349 (L176P_0r, L176P_0a);
  tkr_ra_monitor #("Poly_eval.L176.A") I350 (L176A_0r, L176A_0a);
  tkr_ra_monitor #("Poly_eval.L177.P") I351 (L177P_0r, L177P_0a);
  tkr_ra_monitor #("Poly_eval.L177.A") I352 (L177A_0r, L177A_0a);
  tkr_dr_monitor #("Poly_eval.L178.P", 32) I353 (L178P_0r0[31:0], L178P_0r1[31:0], L178P_0a);
  tkr_dr_monitor #("Poly_eval.L178.A", 32) I354 (L178A_0r0[31:0], L178A_0r1[31:0], L178A_0a);
  tkr_ra_monitor #("Poly_eval.L179.L") I355 (L179_0r, L179_0a);
  tkr_dr_monitor #("Poly_eval.L180.P", 32) I356 (L180P_0r0[31:0], L180P_0r1[31:0], L180P_0a);
  tkr_dr_monitor #("Poly_eval.L180.A", 32) I357 (L180A_0r0[31:0], L180A_0r1[31:0], L180A_0a);
  tkr_dr_monitor #("Poly_eval.L181.P", 2) I358 (L181P_0r0[1:0], L181P_0r1[1:0], L181P_0a);
  tkr_dr_monitor #("Poly_eval.L181.A", 2) I359 (L181A_0r0[1:0], L181A_0r1[1:0], L181A_0a);
  tkr_dr_monitor #("Poly_eval.L182.L", 2) I360 (L182_0r0[1:0], L182_0r1[1:0], L182_0a);
  tkr_dr_monitor #("Poly_eval.L183.P", 2) I361 (L183P_0r0[1:0], L183P_0r1[1:0], L183P_0a);
  tkr_dr_monitor #("Poly_eval.L183.A", 2) I362 (L183A_0r0[1:0], L183A_0r1[1:0], L183A_0a);
  tkr_dr_monitor #("Poly_eval.L184.P", 2) I363 (L184P_0r0[1:0], L184P_0r1[1:0], L184P_0a);
  tkr_dr_monitor #("Poly_eval.L184.A", 2) I364 (L184A_0r0[1:0], L184A_0r1[1:0], L184A_0a);
  tkr_dr_monitor #("Poly_eval.L185.P", 32) I365 (L185P_0r0[31:0], L185P_0r1[31:0], L185P_0a);
  tkr_dr_monitor #("Poly_eval.L185.A", 32) I366 (L185A_0r0[31:0], L185A_0r1[31:0], L185A_0a);
  tkr_ra_monitor #("Poly_eval.L186.P") I367 (L186P_0r, L186P_0a);
  tkr_ra_monitor #("Poly_eval.L186.A") I368 (L186A_0r, L186A_0a);
  tkr_ra_monitor #("Poly_eval.L187.P") I369 (L187P_0r, L187P_0a);
  tkr_ra_monitor #("Poly_eval.L187.A") I370 (L187A_0r, L187A_0a);
  tkr_dr_monitor #("Poly_eval.L188.P", 32) I371 (L188P_0r0[31:0], L188P_0r1[31:0], L188P_0a);
  tkr_dr_monitor #("Poly_eval.L188.A", 32) I372 (L188A_0r0[31:0], L188A_0r1[31:0], L188A_0a);
  tkr_ra_monitor #("Poly_eval.L189.P") I373 (L189P_0r, L189P_0a);
  tkr_ra_monitor #("Poly_eval.L189.A") I374 (L189A_0r, L189A_0a);
  tkr_dr_monitor #("Poly_eval.L190.L", 32) I375 (L190_0r0[31:0], L190_0r1[31:0], L190_0a);
  tkr_ra_monitor #("Poly_eval.L191.L") I376 (L191_0r, L191_0a);
  tkr_dr_monitor #("Poly_eval.L192.L", 32) I377 (L192_0r0[31:0], L192_0r1[31:0], L192_0a);
  tkr_dr_monitor #("Poly_eval.L193.P", 3) I378 (L193P_0r0[2:0], L193P_0r1[2:0], L193P_0a);
  tkr_dr_monitor #("Poly_eval.L193.A", 3) I379 (L193A_0r0[2:0], L193A_0r1[2:0], L193A_0a);
  tkr_dr_monitor #("Poly_eval.L194.P", 3) I380 (L194P_0r0[2:0], L194P_0r1[2:0], L194P_0a);
  tkr_dr_monitor #("Poly_eval.L194.A", 3) I381 (L194A_0r0[2:0], L194A_0r1[2:0], L194A_0a);
  tkr_dr_monitor #("Poly_eval.L195.L", 3) I382 (L195_0r0[2:0], L195_0r1[2:0], L195_0a);
  tkr_dr_monitor #("Poly_eval.L196.P", 3) I383 (L196P_0r0[2:0], L196P_0r1[2:0], L196P_0a);
  tkr_dr_monitor #("Poly_eval.L196.A", 3) I384 (L196A_0r0[2:0], L196A_0r1[2:0], L196A_0a);
  tkr_dr_monitor #("Poly_eval.L197.P", 3) I385 (L197P_0r0[2:0], L197P_0r1[2:0], L197P_0a);
  tkr_dr_monitor #("Poly_eval.L197.A", 3) I386 (L197A_0r0[2:0], L197A_0r1[2:0], L197A_0a);
  tkr_ra_monitor #("Poly_eval.L198.P") I387 (L198P_0r, L198P_0a);
  tkr_ra_monitor #("Poly_eval.L198.A") I388 (L198A_0r, L198A_0a);
  tkr_dr_monitor #("Poly_eval.L199.L", 32) I389 (L199_0r0[31:0], L199_0r1[31:0], L199_0a);
  tkr_ra_monitor #("Poly_eval.L200.L") I390 (L200_0r, L200_0a);
  tkr_dr_monitor #("Poly_eval.L206.L", 64) I391 (L206_0r0[63:0], L206_0r1[63:0], L206_0a);
  tkr_dr_monitor #("Poly_eval.L211.L", 32) I392 (L211_0r0[31:0], L211_0r1[31:0], L211_0a);
  tkr_ra_monitor #("Poly_eval.L216.L") I393 (L216_0r, L216_0a);
  tkr_ra_monitor #("Poly_eval.L217.L") I394 (L217_0r, L217_0a);
  tkr_ra_monitor #("Poly_eval.L218.L") I395 (L218_0r, L218_0a);
  tkr_dr_monitor #("Poly_eval.L224.L", 64) I396 (L224_0r0[63:0], L224_0r1[63:0], L224_0a);
  tkr_dr_monitor #("Poly_eval.L229.L", 32) I397 (L229_0r0[31:0], L229_0r1[31:0], L229_0a);
  tkr_ra_monitor #("Poly_eval.L234.L") I398 (L234_0r, L234_0a);
  tkr_ra_monitor #("Poly_eval.L235.L") I399 (L235_0r, L235_0a);
  tkr_ra_monitor #("Poly_eval.L236.L") I400 (L236_0r, L236_0a);
  tkr_dr_monitor #("Poly_eval.L242.L", 64) I401 (L242_0r0[63:0], L242_0r1[63:0], L242_0a);
  tkr_dr_monitor #("Poly_eval.L247.L", 32) I402 (L247_0r0[31:0], L247_0r1[31:0], L247_0a);
  tkr_dr_monitor #("Poly_eval.L249.L", 32) I403 (L249_0r0[31:0], L249_0r1[31:0], L249_0a);
  tkr_ra_monitor #("Poly_eval.L252.L") I404 (L252_0r, L252_0a);
  tkr_ra_monitor #("Poly_eval.L253.P") I405 (L253P_0r, L253P_0a);
  tkr_ra_monitor #("Poly_eval.L253.A") I406 (L253A_0r, L253A_0a);
  tkr_ra_monitor #("Poly_eval.L254.L") I407 (L254_0r, L254_0a);
  tkr_ra_monitor #("Poly_eval.L255.P") I408 (L255P_0r, L255P_0a);
  tkr_ra_monitor #("Poly_eval.L255.A") I409 (L255A_0r, L255A_0a);
  tkr_ra_monitor #("Poly_eval.L257.P") I410 (L257P_0r, L257P_0a);
  tkr_ra_monitor #("Poly_eval.L257.A") I411 (L257A_0r, L257A_0a);
  tkr_ra_monitor #("Poly_eval.L260.P") I412 (L260P_0r, L260P_0a);
  tkr_ra_monitor #("Poly_eval.L260.A") I413 (L260A_0r, L260A_0a);
  tkr_dr_monitor #("Poly_eval.L264.P", 32) I414 (L264P_0r0[31:0], L264P_0r1[31:0], L264P_0a);
  tkr_dr_monitor #("Poly_eval.L264.A", 32) I415 (L264A_0r0[31:0], L264A_0r1[31:0], L264A_0a);
  tkr_ra_monitor #("Poly_eval.L267.L") I416 (L267_0r, L267_0a);
  tkr_dr_monitor #("Poly_eval.L272.P", 33) I417 (L272P_0r0[32:0], L272P_0r1[32:0], L272P_0a);
  tkr_dr_monitor #("Poly_eval.L272.A", 33) I418 (L272A_0r0[32:0], L272A_0r1[32:0], L272A_0a);
  tkr_ra_monitor #("Poly_eval.L275.P") I419 (L275P_0r, L275P_0a);
  tkr_ra_monitor #("Poly_eval.L275.A") I420 (L275A_0r, L275A_0a);
  tkr_ra_monitor #("Poly_eval.L277.P") I421 (L277P_0r, L277P_0a);
  tkr_ra_monitor #("Poly_eval.L277.A") I422 (L277A_0r, L277A_0a);
  tkr_ra_monitor #("Poly_eval.L278.L") I423 (L278_0r, L278_0a);
  tkr_ra_monitor #("Poly_eval.L281.P") I424 (L281P_0r, L281P_0a);
  tkr_ra_monitor #("Poly_eval.L281.A") I425 (L281A_0r, L281A_0a);
  tkr_ra_monitor #("Poly_eval.L284.P") I426 (L284P_0r, L284P_0a);
  tkr_ra_monitor #("Poly_eval.L284.A") I427 (L284A_0r, L284A_0a);
  tkr_dr_monitor #("Poly_eval.L286.L", 32) I428 (L286_0r0[31:0], L286_0r1[31:0], L286_0a);
  tkr_dr_monitor #("Poly_eval.L288.L", 32) I429 (L288_0r0[31:0], L288_0r1[31:0], L288_0a);
  tkr_dr_monitor #("Poly_eval.L289.L", 3) I430 (L289_0r0[2:0], L289_0r1[2:0], L289_0a);
  tkr_dr_monitor #("Poly_eval.L290.L", 3) I431 (L290_0r0[2:0], L290_0r1[2:0], L290_0a);
  tkr_dr_monitor #("Poly_eval.L291.L", 3) I432 (L291_0r0[2:0], L291_0r1[2:0], L291_0a);
  tkr_dr_monitor #("Poly_eval.L292.L", 3) I433 (L292_0r0[2:0], L292_0r1[2:0], L292_0a);
  tkr_dr_monitor #("Poly_eval.L293.L", 35) I434 (L293_0r0[34:0], L293_0r1[34:0], L293_0a);
  tkr_dr_monitor #("Poly_eval.L295.L", 32) I435 (L295_0r0[31:0], L295_0r1[31:0], L295_0a);
  tkr_dr_monitor #("Poly_eval.L297.L", 32) I436 (L297_0r0[31:0], L297_0r1[31:0], L297_0a);
  tkr_dr_monitor #("Poly_eval.L299.L", 32) I437 (L299_0r0[31:0], L299_0r1[31:0], L299_0a);
  tkr_dr_monitor #("Poly_eval.L302.P", 32) I438 (L302P_0r0[31:0], L302P_0r1[31:0], L302P_0a);
  tkr_dr_monitor #("Poly_eval.L302.A", 32) I439 (L302A_0r0[31:0], L302A_0r1[31:0], L302A_0a);
  tkr_dr_monitor #("Poly_eval.L308.P", 32) I440 (L308P_0r0[31:0], L308P_0r1[31:0], L308P_0a);
  tkr_dr_monitor #("Poly_eval.L308.A", 32) I441 (L308A_0r0[31:0], L308A_0r1[31:0], L308A_0a);
  tkr_ra_monitor #("Poly_eval.L309.L") I442 (L309_0r, L309_0a);
  tkr_ra_monitor #("Poly_eval.L310.L") I443 (L310_0r, L310_0a);
  tkr_dr_monitor #("Poly_eval.L311.L", 32) I444 (L311_0r0[31:0], L311_0r1[31:0], L311_0a);
  tkr_ra_monitor #("Poly_eval.L312.L") I445 (L312_0r, L312_0a);
  tkr_dr_monitor #("Poly_eval.L313.P", 32) I446 (L313P_0r0[31:0], L313P_0r1[31:0], L313P_0a);
  tkr_dr_monitor #("Poly_eval.L313.A", 32) I447 (L313A_0r0[31:0], L313A_0r1[31:0], L313A_0a);
  tkr_dr_monitor #("Poly_eval.L314.L", 2) I448 (L314_0r0[1:0], L314_0r1[1:0], L314_0a);
  tkr_dr_monitor #("Poly_eval.L315.L", 2) I449 (L315_0r0[1:0], L315_0r1[1:0], L315_0a);
  tkr_dr_monitor #("Poly_eval.L316.L", 2) I450 (L316_0r0[1:0], L316_0r1[1:0], L316_0a);
  tkr_dr_monitor #("Poly_eval.L317.P", 2) I451 (L317P_0r0[1:0], L317P_0r1[1:0], L317P_0a);
  tkr_dr_monitor #("Poly_eval.L317.A", 2) I452 (L317A_0r0[1:0], L317A_0r1[1:0], L317A_0a);
  tkr_dr_monitor #("Poly_eval.L318.P", 32) I453 (L318P_0r0[31:0], L318P_0r1[31:0], L318P_0a);
  tkr_dr_monitor #("Poly_eval.L318.A", 32) I454 (L318A_0r0[31:0], L318A_0r1[31:0], L318A_0a);
  tkr_ra_monitor #("Poly_eval.L319.P") I455 (L319P_0r, L319P_0a);
  tkr_ra_monitor #("Poly_eval.L319.A") I456 (L319A_0r, L319A_0a);
  tkr_ra_monitor #("Poly_eval.L320.P") I457 (L320P_0r, L320P_0a);
  tkr_ra_monitor #("Poly_eval.L320.A") I458 (L320A_0r, L320A_0a);
  tkr_dr_monitor #("Poly_eval.L321.L", 32) I459 (L321_0r0[31:0], L321_0r1[31:0], L321_0a);
  tkr_ra_monitor #("Poly_eval.L322.L") I460 (L322_0r, L322_0a);
  tkr_dr_monitor #("Poly_eval.L323.L", 32) I461 (L323_0r0[31:0], L323_0r1[31:0], L323_0a);
  tkr_dr_monitor #("Poly_eval.L324.P", 2) I462 (L324P_0r0[1:0], L324P_0r1[1:0], L324P_0a);
  tkr_dr_monitor #("Poly_eval.L324.A", 2) I463 (L324A_0r0[1:0], L324A_0r1[1:0], L324A_0a);
  tkr_dr_monitor #("Poly_eval.L325.L", 2) I464 (L325_0r0[1:0], L325_0r1[1:0], L325_0a);
  tkr_dr_monitor #("Poly_eval.L326.P", 2) I465 (L326P_0r0[1:0], L326P_0r1[1:0], L326P_0a);
  tkr_dr_monitor #("Poly_eval.L326.A", 2) I466 (L326A_0r0[1:0], L326A_0r1[1:0], L326A_0a);
  tkr_dr_monitor #("Poly_eval.L327.P", 2) I467 (L327P_0r0[1:0], L327P_0r1[1:0], L327P_0a);
  tkr_dr_monitor #("Poly_eval.L327.A", 2) I468 (L327A_0r0[1:0], L327A_0r1[1:0], L327A_0a);
  tkr_dr_monitor #("Poly_eval.L328.L", 32) I469 (x_0r0[31:0], x_0r1[31:0], x_0a);
  tkr_dr_monitor #("Poly_eval.L329.L", 32) I470 (coefs_0_0r0[31:0], coefs_0_0r1[31:0], coefs_0_0a);
  tkr_dr_monitor #("Poly_eval.L330.L", 32) I471 (coefs_1_0r0[31:0], coefs_1_0r1[31:0], coefs_1_0a);
  tkr_dr_monitor #("Poly_eval.L331.L", 32) I472 (coefs_2_0r0[31:0], coefs_2_0r1[31:0], coefs_2_0a);
  tkr_dr_monitor #("Poly_eval.L332.L", 2) I473 (L332_0r0[1:0], L332_0r1[1:0], L332_0a);
  tkr_dr_monitor #("Poly_eval.L333.P", 2) I474 (L333P_0r0[1:0], L333P_0r1[1:0], L333P_0a);
  tkr_dr_monitor #("Poly_eval.L333.A", 2) I475 (L333A_0r0[1:0], L333A_0r1[1:0], L333A_0a);
  tkr_dr_monitor #("Poly_eval.L334.P", 2) I476 (L334P_0r0[1:0], L334P_0r1[1:0], L334P_0a);
  tkr_dr_monitor #("Poly_eval.L334.A", 2) I477 (L334A_0r0[1:0], L334A_0r1[1:0], L334A_0a);
  tkr_dr_monitor #("Poly_eval.L335.L", 34) I478 (L335_0r0[33:0], L335_0r1[33:0], L335_0a);
  tkr_dr_monitor #("Poly_eval.L336.L", 32) I479 (a_0r0[31:0], a_0r1[31:0], a_0a);
  tkr_ra_monitor #("Poly_eval.L338.P") I480 (L338P_0r, L338P_0a);
  tkr_ra_monitor #("Poly_eval.L338.A") I481 (L338A_0r, L338A_0a);
  tkr_dr_monitor #("Poly_eval.L345.P", 1) I482 (L345P_0r0, L345P_0r1, L345P_0a);
  tkr_dr_monitor #("Poly_eval.L345.A", 1) I483 (L345A_0r0, L345A_0r1, L345A_0a);
  tkr_dr_monitor #("Poly_eval.L346.P", 1) I484 (L346P_0r0, L346P_0r1, L346P_0a);
  tkr_dr_monitor #("Poly_eval.L346.A", 1) I485 (L346A_0r0, L346A_0r1, L346A_0a);
  tkr_dr_monitor #("Poly_eval.L347.P", 3) I486 (L347P_0r0[2:0], L347P_0r1[2:0], L347P_0a);
  tkr_dr_monitor #("Poly_eval.L347.A", 3) I487 (L347A_0r0[2:0], L347A_0r1[2:0], L347A_0a);
  tkr_dr_monitor #("Poly_eval.L348.P", 1) I488 (L348P_0r0, L348P_0r1, L348P_0a);
  tkr_dr_monitor #("Poly_eval.L348.A", 1) I489 (L348A_0r0, L348A_0r1, L348A_0a);
  tkr_dr_monitor #("Poly_eval.L349.L", 3) I490 (L349_0r0[2:0], L349_0r1[2:0], L349_0a);
  tkr_dr_monitor #("Poly_eval.L350.L", 32) I491 (L350_0r0[31:0], L350_0r1[31:0], L350_0a);
  tkr_dr_monitor #("Poly_eval.L351.L", 32) I492 (L351_0r0[31:0], L351_0r1[31:0], L351_0a);
  tkr_dr_monitor #("Poly_eval.L352.L", 3) I493 (L352_0r0[2:0], L352_0r1[2:0], L352_0a);
  tkr_dr_monitor #("Poly_eval.L353.P", 32) I494 (L353P_0r0[31:0], L353P_0r1[31:0], L353P_0a);
  tkr_dr_monitor #("Poly_eval.L353.A", 32) I495 (L353A_0r0[31:0], L353A_0r1[31:0], L353A_0a);
  tkr_ra_monitor #("Poly_eval.L355.L") I496 (L355_0r, L355_0a);
  tkr_ra_monitor #("Poly_eval.L356.L") I497 (L356_0r, L356_0a);
  tkr_ra_monitor #("Poly_eval.L357.L") I498 (L357_0r, L357_0a);
  tkr_dr_monitor #("Poly_eval.L358.P", 32) I499 (L358P_0r0[31:0], L358P_0r1[31:0], L358P_0a);
  tkr_dr_monitor #("Poly_eval.L358.A", 32) I500 (L358A_0r0[31:0], L358A_0r1[31:0], L358A_0a);
  tkr_dr_monitor #("Poly_eval.L359.P", 32) I501 (L359P_0r0[31:0], L359P_0r1[31:0], L359P_0a);
  tkr_dr_monitor #("Poly_eval.L359.A", 32) I502 (L359A_0r0[31:0], L359A_0r1[31:0], L359A_0a);
  tkr_dr_monitor #("Poly_eval.L360.P", 32) I503 (L360P_0r0[31:0], L360P_0r1[31:0], L360P_0a);
  tkr_dr_monitor #("Poly_eval.L360.A", 32) I504 (L360A_0r0[31:0], L360A_0r1[31:0], L360A_0a);
  tkr_ra_monitor #("Poly_eval.L361.P") I505 (L361P_0r, L361P_0a);
  tkr_ra_monitor #("Poly_eval.L361.A") I506 (L361A_0r, L361A_0a);
  tkr_ra_monitor #("Poly_eval.L362.P") I507 (L362P_0r, L362P_0a);
  tkr_ra_monitor #("Poly_eval.L362.A") I508 (L362A_0r, L362A_0a);
  tkr_ra_monitor #("Poly_eval.L363.P") I509 (L363P_0r, L363P_0a);
  tkr_ra_monitor #("Poly_eval.L363.A") I510 (L363A_0r, L363A_0a);
  tkr_ra_monitor #("Poly_eval.L364.P") I511 (L364P_0r, L364P_0a);
  tkr_ra_monitor #("Poly_eval.L364.A") I512 (L364A_0r, L364A_0a);
  tkr_ra_monitor #("Poly_eval.L366.P") I513 (L366P_0r, L366P_0a);
  tkr_ra_monitor #("Poly_eval.L366.A") I514 (L366A_0r, L366A_0a);
  tkr_ra_monitor #("Poly_eval.L367.P") I515 (L367P_0r, L367P_0a);
  tkr_ra_monitor #("Poly_eval.L367.A") I516 (L367A_0r, L367A_0a);
  tkr_ra_monitor #("Poly_eval.L385.P") I517 (L385P_0r, L385P_0a);
  tkr_ra_monitor #("Poly_eval.L385.A") I518 (L385A_0r, L385A_0a);
  tkr_dr_monitor #("Poly_eval.L395.P", 32) I519 (L395P_0r0[31:0], L395P_0r1[31:0], L395P_0a);
  tkr_dr_monitor #("Poly_eval.L395.A", 32) I520 (L395A_0r0[31:0], L395A_0r1[31:0], L395A_0a);
endmodule

// Netlist costs:
// teak_Poly_eval: AND2*2914 AO22*205 AO222*582 BUFF*4413 C2*1035 C2R*1846 C3*3983 GND*329 INV*701 NAND2*588 NAND3*12 NOR2*224 NOR3*822 OR2*2289 OR3*248
// tkf0mo0w0_o0w0: BUFF*2 C2*1
// tkf0mo0w0_o0w0_o0w0: BUFF*3 C3*1
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0: BUFF*5 C2*2 C3*1
// tkf32mo0w0_o0w32: BUFF*66 C3*1 OR2*1
// tkf33mo0w0_o0w32: BUFF*64 C2*3 C3*1 OR2*2
// tkf4mo0w0_o0w3: BUFF*6 C2*3 C3*1 OR2*2
// tki: AND2*1 AO22*3 INV*3
// tkj0m0_0: BUFF*2 C2*1
// tkj2m0_2: BUFF*9 C2*2
// tkj32m32_0: BUFF*129 C2*2
// tkj32m32_0_0_0: BUFF*130 C2*2 C3*1
// tkj34m32_2: BUFF*137 C2*2 OR2*1
// tkj35m32_3: BUFF*141 C2*2 OR2*1
// tkj3m0_3: BUFF*13 C2*2
// tkj64m32_32: BUFF*257 C2*2 OR2*1
// tkj64m32_32_0: BUFF*257 C2*3 OR2*1
// tkl0x1: BUFF*1 C2R*1 INV*1
// tkl1x1: BUFF*1 C2R*2 INV*1 OR2*1
// tkl2x1: C2*1 C2R*4 INV*1 OR2*2
// tkl32x1: BUFF*1 C2*3 C2R*64 C3*14 INV*1 OR2*32
// tkl33x1: BUFF*1 C2*2 C2R*66 C3*15 INV*1 OR2*33
// tkl3x1: C2R*6 C3*1 INV*1 OR2*3
// tkl4x1: BUFF*1 C2*1 C2R*8 C3*1 INV*1 OR2*4
// tkl64x1: BUFF*2 C2*1 C2R*128 C3*31 INV*1 OR2*64
// tkm2x0b: C2R*4 NOR2*1 OR2*1
// tkm2x2b: AND2*8 C2*2 C2R*4 NOR2*1 OR2*9
// tkm2x32b: AND2*128 BUFF*2 C2*6 C2R*4 C3*28 NOR2*1 OR2*129
// tkm3x0b: C2R*6 NOR2*1 OR3*1
// tkm3x32b: AND2*192 BUFF*3 C2*9 C2R*6 C3*42 NOR2*1 OR2*96 OR3*65
// tkm3x3b: AND2*18 C2R*6 C3*3 NOR2*1 OR2*9 OR3*7
// tko0m2_1nm2b1: BUFF*3 GND*2
// tko0m2_1nm2b2: BUFF*3 GND*2
// tko0m32_1nm32b0: BUFF*33 GND*32
// tko0m32_1nm32b1: BUFF*33 GND*32
// tko0m3_1nm3b0: BUFF*4 GND*3
// tko0m3_1nm3b1: BUFF*4 GND*3
// tko0m3_1nm3b2: BUFF*4 GND*3
// tko0m3_1nm3b4: BUFF*4 GND*3
// tko1m1_1nm1b1_2eqi0w1bt1o0w1b: BUFF*5 C2*4 GND*1 OR2*3
// tko1m1_1nm1b1_2nei0w1bt1o0w1b: BUFF*5 C2*4 GND*1 OR2*3
// tko32m1_1nm32b0_2sgti0w32bt1o0w32b: BUFF*35 C2*224 C3*14 GND*32 OR2*127
// tko32m32_1nm32b0_2subt1o0w32bi0w32b: AO222*62 BUFF*35 C2*7 C3*262 GND*32 INV*62 NAND2*62 NOR3*62 OR2*34 OR3*1
// tko32m33_1api0w32bi31w1b_2nm33b1_3subt1o0w33bt2o0w33b: AO222*64 BUFF*102 C2*7 C3*270 GND*33 INV*64 NAND2*64 NOR3*64 OR2*34 OR3*1
// tko3m1_1nm3b1_2eqi0w3bt1o0w3b: BUFF*8 C2*20 C3*1 GND*3 OR2*9 OR3*2
// tko3m4_1nm1b0_2api0w3bt1o0w1b_3nm4b1_4addt2o0w4bt3o0w4b: AO222*6 BUFF*15 C2*4 C3*25 GND*5 INV*6 NAND2*6 NOR3*6 OR2*5 OR3*1
// tko64m32_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b_4apt3o0w32b: AO222*64 BUFF*198 C2*4 C3*256 INV*64 NAND2*64 NOR3*64 OR2*2 OR3*1
// tko64m33_1api0w32bi31w1b_2api32w32bi63w1b_3addt1o0w33bt2o0w33b: AO222*64 BUFF*134 C2*4 C3*256 INV*64 NAND2*64 NOR3*64 OR2*2 OR3*1
// tks1_o0w1_0o0w0_1o0w0: BUFF*7 C2*3 OR2*2
// tks2_o0w2_1o0w0_2o0w0: BUFF*4 C2*6 OR2*3
// tks32_o0w32_3cfffffffcm4cfffffff8m5cfffffff8m6cfffffff8m8cfffffff0m9cfffffff0macfffffff0m10cffffffe0m11cffffffe0m12cffffffe0m20cffffffc0m21cffffffc0m22cffffffc0m40cffffff80m41cffffff80m42cffffff80m80cffffff00m81cffffff00m82cffffff00m100cfffffe00m101cfffffe00m102cfffffe00m200cfffffc00m201cfffffc00m202cfffffc00m400cfffff800m401cfffff800m402cfffff800m800cfffff000m801cfffff000m802cfffff000m1000cffffe000m1001cffffe000m1002cffffe000m2000cffffc000m2001cffffc000m2002cffffc000m4000cffff8000m4001cffff8000m4002cffff8000m8000cffff0000m8001cffff0000m8002cffff0000m10000cfffe0000m10001cfffe0000m10002cfffe0000m20000cfffc0000m20001cfffc0000m20002cfffc0000m40000cfff80000m40001cfff80000m40002cfff80000m80000cfff00000m80001cfff00000m80002cfff00000m100000cffe00000m100001cffe00000m100002cffe00000m200000cffc00000m200001cffc00000m200002cffc00000m400000cff800000m400001cff800000m400002cff800000m800000cff000000m800001cff000000m800002cff000000m1000000cfe000000m1000001cfe000000m1000002cfe000000m2000000cfc000000m2000001cfc000000m2000002cfc000000m4000000cf8000000m4000001cf8000000m4000002cf8000000m8000000cf0000000m8000001cf0000000m8000002cf0000000m10000000ce0000000m10000001ce0000000m10000002ce0000000m20000000cc0000000m20000001cc0000000m20000002cc0000000m40000000c80000000m40000001c80000000m40000002c80000000m80000000m80000001m80000002o0w0_0o0w0_1o0w0_2o0w0: BUFF*83 C2*123 C3*746 INV*4 NAND2*1 NAND3*11 NOR2*1 NOR3*34 OR2*33
// tks34_o32w2_1o0w32_2o0w32: BUFF*4 C2*134 C3*16 OR2*35
// tks35_o32w3_1o0w32_2o0w32_4o0w32: BUFF*4 C2*198 C3*19 OR2*35 OR3*1
// tks3_o0w3_1o0w0_2o0w0_4o0w0: BUFF*6 C2*4 C3*4 OR2*3 OR3*1
// tkvaV32_wo0w32_ro0w32o0w32: AND2*288 AO22*33 BUFF*102 C2*5 C3*29 INV*2 NAND2*1 NOR2*33 NOR3*33 OR2*32
// tkvi32_wo0w32_ro0w32o0w32o31w1: AND2*290 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvneg3_wo0w3_ro0w3o0w3o0w3: AND2*33 AO22*4 BUFF*15 C2*1 C3*2 INV*1 NAND2*1 NOR2*4 NOR3*5 OR2*3
// tkvr132_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvr232_wo0w32_ro0w32o0w32o31w1: AND2*290 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvr332_wo0w32_ro0w32o0w32o0w32o31w1: AND2*354 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvxV32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
